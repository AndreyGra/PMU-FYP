// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition"

// DATE "03/10/2020 09:20:21"

// 
// Device: Altera 5CSEMA6F31C8 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module IoTOctopus_QSYS (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_32_clk,
	mac_mdio_connection_mdc,
	mac_mdio_connection_mdio_in,
	mac_mdio_connection_mdio_out,
	mac_mdio_connection_mdio_oen,
	mac_misc_connection_magic_wakeup,
	mac_misc_connection_magic_sleep_n,
	mac_misc_connection_ff_tx_crc_fwd,
	mac_misc_connection_ff_tx_septy,
	mac_misc_connection_tx_ff_uflow,
	mac_misc_connection_ff_tx_a_full,
	mac_misc_connection_ff_tx_a_empty,
	mac_misc_connection_rx_err_stat,
	mac_misc_connection_rx_frm_type,
	mac_misc_connection_ff_rx_dsav,
	mac_misc_connection_ff_rx_a_full,
	mac_misc_connection_ff_rx_a_empty,
	mac_rgmii_connection_rgmii_in,
	mac_rgmii_connection_rgmii_out,
	mac_rgmii_connection_rx_control,
	mac_rgmii_connection_tx_control,
	mac_rx_clock_connection_clk,
	mac_status_connection_set_10,
	mac_status_connection_set_1000,
	mac_status_connection_eth_mode,
	mac_status_connection_ena_10,
	mac_tx_clock_connection_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_32_clk;
output 	mac_mdio_connection_mdc;
input 	mac_mdio_connection_mdio_in;
output 	mac_mdio_connection_mdio_out;
output 	mac_mdio_connection_mdio_oen;
output 	mac_misc_connection_magic_wakeup;
input 	mac_misc_connection_magic_sleep_n;
input 	mac_misc_connection_ff_tx_crc_fwd;
output 	mac_misc_connection_ff_tx_septy;
output 	mac_misc_connection_tx_ff_uflow;
output 	mac_misc_connection_ff_tx_a_full;
output 	mac_misc_connection_ff_tx_a_empty;
output 	[17:0] mac_misc_connection_rx_err_stat;
output 	[3:0] mac_misc_connection_rx_frm_type;
output 	mac_misc_connection_ff_rx_dsav;
output 	mac_misc_connection_ff_rx_a_full;
output 	mac_misc_connection_ff_rx_a_empty;
input 	[3:0] mac_rgmii_connection_rgmii_in;
output 	[3:0] mac_rgmii_connection_rgmii_out;
input 	mac_rgmii_connection_rx_control;
output 	mac_rgmii_connection_tx_control;
input 	mac_rx_clock_connection_clk;
input 	mac_status_connection_set_10;
input 	mac_status_connection_set_1000;
output 	mac_status_connection_eth_mode;
output 	mac_status_connection_ena_10;
input 	mac_tx_clock_connection_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[0] ;
wire \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[1] ;
wire \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[2] ;
wire \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[3] ;
wire \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out1|altddio_out_component|auto_generated|dataout[0] ;
wire \eth_tse_0|i_tse_mac|U_MDIO|U_CLKGEN|mdio_clk~q ;
wire \eth_tse_0|i_tse_mac|U_MDIO|mdio_out~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|command_config[21]~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|septy_flag~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_GETH|U_TX|tx_ff_uflow~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|afull_flag~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|aempty_flag~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|state.LOC_STATE_DATA~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|state.LOC_STATE_SHIFT~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[5]~0_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[6]~1_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[7]~2_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[8]~3_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[9]~4_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[10]~5_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[11]~6_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[12]~7_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[13]~8_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[14]~9_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[15]~10_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[16]~11_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[17]~12_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[18]~13_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[19]~14_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[20]~15_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[4]~16_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[22]~17_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_ucast~0_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_mcast~0_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_bcast~0_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_vlan~0_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|sav_flag~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|afull_flag~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|aempty_flag~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|eth_mode~q ;
wire \eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|ena_10~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \avalon_st_adapter_001|timing_adapter_0|LessThan0~0_combout ;
wire \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|U_SYNC_2|sync[10].u|std_sync_no_cut|din_s1~0_combout ;
wire \~GND~combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \mac_mdio_connection_mdio_in~input_o ;
wire \clk_32_clk~input_o ;
wire \mac_tx_clock_connection_clk~input_o ;
wire \mac_rx_clock_connection_clk~input_o ;
wire \mac_status_connection_set_1000~input_o ;
wire \mac_status_connection_set_10~input_o ;
wire \reset_reset_n~input_o ;
wire \mac_misc_connection_ff_tx_crc_fwd~input_o ;
wire \mac_rgmii_connection_rgmii_in[3]~input_o ;
wire \mac_rgmii_connection_rgmii_in[2]~input_o ;
wire \mac_rgmii_connection_rgmii_in[1]~input_o ;
wire \mac_rgmii_connection_rgmii_in[0]~input_o ;
wire \mac_rgmii_connection_rx_control~input_o ;
wire \mac_misc_connection_magic_sleep_n~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|BWHK8171_1~q ;
wire \nabboc|pzdyqx_impl_inst|BWHK8171_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ZIVV0726~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ZIVV0726~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12_combout ;
wire \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ;
wire \nabboc|pzdyqx_impl_inst|sdr~combout ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1]~q ;
wire \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


IoTOctopus_QSYS_altera_reset_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_32_clk(\clk_32_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

IoTOctopus_QSYS_IoTOctopus_QSYS_avalon_st_adapter_001 avalon_st_adapter_001(
	.stateLOC_STATE_DATA(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|state.LOC_STATE_DATA~q ),
	.stateLOC_STATE_SHIFT(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|state.LOC_STATE_SHIFT~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.LessThan0(\avalon_st_adapter_001|timing_adapter_0|LessThan0~0_combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk_32_clk(\clk_32_clk~input_o ));

IoTOctopus_QSYS_IoTOctopus_QSYS_eth_tse_0 eth_tse_0(
	.dataout_0(\eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[0] ),
	.dataout_1(\eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[1] ),
	.dataout_2(\eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[2] ),
	.dataout_3(\eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[3] ),
	.dataout_01(\eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out1|altddio_out_component|auto_generated|dataout[0] ),
	.mdio_clk(\eth_tse_0|i_tse_mac|U_MDIO|U_CLKGEN|mdio_clk~q ),
	.mdio_out(\eth_tse_0|i_tse_mac|U_MDIO|mdio_out~q ),
	.command_config_21(\eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|command_config[21]~q ),
	.septy_flag(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|septy_flag~q ),
	.tx_ff_uflow(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_GETH|U_TX|tx_ff_uflow~q ),
	.afull_flag(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|afull_flag~q ),
	.aempty_flag(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|aempty_flag~q ),
	.stateLOC_STATE_DATA(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|state.LOC_STATE_DATA~q ),
	.stateLOC_STATE_SHIFT(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|state.LOC_STATE_SHIFT~q ),
	.ff_rx_err_stat_5(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[5]~0_combout ),
	.ff_rx_err_stat_6(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[6]~1_combout ),
	.ff_rx_err_stat_7(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[7]~2_combout ),
	.ff_rx_err_stat_8(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[8]~3_combout ),
	.ff_rx_err_stat_9(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[9]~4_combout ),
	.ff_rx_err_stat_10(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[10]~5_combout ),
	.ff_rx_err_stat_11(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[11]~6_combout ),
	.ff_rx_err_stat_12(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[12]~7_combout ),
	.ff_rx_err_stat_13(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[13]~8_combout ),
	.ff_rx_err_stat_14(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[14]~9_combout ),
	.ff_rx_err_stat_15(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[15]~10_combout ),
	.ff_rx_err_stat_16(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[16]~11_combout ),
	.ff_rx_err_stat_17(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[17]~12_combout ),
	.ff_rx_err_stat_18(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[18]~13_combout ),
	.ff_rx_err_stat_19(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[19]~14_combout ),
	.ff_rx_err_stat_20(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[20]~15_combout ),
	.ff_rx_err_stat_4(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[4]~16_combout ),
	.ff_rx_err_stat_22(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[22]~17_combout ),
	.ff_rx_ucast(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_ucast~0_combout ),
	.ff_rx_mcast(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_mcast~0_combout ),
	.ff_rx_bcast(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_bcast~0_combout ),
	.ff_rx_vlan(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_vlan~0_combout ),
	.sav_flag(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|sav_flag~q ),
	.afull_flag1(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|afull_flag~q ),
	.aempty_flag1(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|aempty_flag~q ),
	.eth_mode(\eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|eth_mode~q ),
	.ena_10(\eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|ena_10~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.LessThan0(\avalon_st_adapter_001|timing_adapter_0|LessThan0~0_combout ),
	.din_s1(\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|U_SYNC_2|sync[10].u|std_sync_no_cut|din_s1~0_combout ),
	.GND_port(\~GND~combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.clk_32_clk(\clk_32_clk~input_o ),
	.mac_tx_clock_connection_clk(\mac_tx_clock_connection_clk~input_o ),
	.mac_rx_clock_connection_clk(\mac_rx_clock_connection_clk~input_o ),
	.mac_status_connection_set_1000(\mac_status_connection_set_1000~input_o ),
	.mac_status_connection_set_10(\mac_status_connection_set_10~input_o ),
	.mac_misc_connection_ff_tx_crc_fwd(\mac_misc_connection_ff_tx_crc_fwd~input_o ),
	.mac_rgmii_connection_rgmii_in_3(\mac_rgmii_connection_rgmii_in[3]~input_o ),
	.mac_rgmii_connection_rgmii_in_2(\mac_rgmii_connection_rgmii_in[2]~input_o ),
	.mac_rgmii_connection_rgmii_in_1(\mac_rgmii_connection_rgmii_in[1]~input_o ),
	.mac_rgmii_connection_rgmii_in_0(\mac_rgmii_connection_rgmii_in[0]~input_o ),
	.mac_rgmii_connection_rx_control(\mac_rgmii_connection_rx_control~input_o ),
	.mac_misc_connection_magic_sleep_n(\mac_misc_connection_magic_sleep_n~input_o ));

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

assign \clk_32_clk~input_o  = clk_32_clk;

assign \mac_tx_clock_connection_clk~input_o  = mac_tx_clock_connection_clk;

assign \mac_rx_clock_connection_clk~input_o  = mac_rx_clock_connection_clk;

assign \mac_status_connection_set_1000~input_o  = mac_status_connection_set_1000;

assign \mac_status_connection_set_10~input_o  = mac_status_connection_set_10;

assign \reset_reset_n~input_o  = reset_reset_n;

assign \mac_misc_connection_ff_tx_crc_fwd~input_o  = mac_misc_connection_ff_tx_crc_fwd;

assign \mac_rgmii_connection_rgmii_in[3]~input_o  = mac_rgmii_connection_rgmii_in[3];

assign \mac_rgmii_connection_rgmii_in[2]~input_o  = mac_rgmii_connection_rgmii_in[2];

assign \mac_rgmii_connection_rgmii_in[1]~input_o  = mac_rgmii_connection_rgmii_in[1];

assign \mac_rgmii_connection_rgmii_in[0]~input_o  = mac_rgmii_connection_rgmii_in[0];

assign \mac_rgmii_connection_rx_control~input_o  = mac_rgmii_connection_rx_control;

assign \mac_misc_connection_magic_sleep_n~input_o  = mac_misc_connection_magic_sleep_n;

assign mac_mdio_connection_mdc = \eth_tse_0|i_tse_mac|U_MDIO|U_CLKGEN|mdio_clk~q ;

assign mac_mdio_connection_mdio_out = \eth_tse_0|i_tse_mac|U_MDIO|mdio_out~q ;

assign mac_mdio_connection_mdio_oen = vcc;

assign mac_misc_connection_magic_wakeup = \eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|command_config[21]~q ;

assign mac_misc_connection_ff_tx_septy = ~ \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|septy_flag~q ;

assign mac_misc_connection_tx_ff_uflow = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_GETH|U_TX|tx_ff_uflow~q ;

assign mac_misc_connection_ff_tx_a_full = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|afull_flag~q ;

assign mac_misc_connection_ff_tx_a_empty = ~ \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|TX_DATA|aempty_flag~q ;

assign mac_misc_connection_rx_err_stat[0] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[5]~0_combout ;

assign mac_misc_connection_rx_err_stat[1] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[6]~1_combout ;

assign mac_misc_connection_rx_err_stat[2] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[7]~2_combout ;

assign mac_misc_connection_rx_err_stat[3] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[8]~3_combout ;

assign mac_misc_connection_rx_err_stat[4] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[9]~4_combout ;

assign mac_misc_connection_rx_err_stat[5] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[10]~5_combout ;

assign mac_misc_connection_rx_err_stat[6] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[11]~6_combout ;

assign mac_misc_connection_rx_err_stat[7] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[12]~7_combout ;

assign mac_misc_connection_rx_err_stat[8] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[13]~8_combout ;

assign mac_misc_connection_rx_err_stat[9] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[14]~9_combout ;

assign mac_misc_connection_rx_err_stat[10] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[15]~10_combout ;

assign mac_misc_connection_rx_err_stat[11] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[16]~11_combout ;

assign mac_misc_connection_rx_err_stat[12] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[17]~12_combout ;

assign mac_misc_connection_rx_err_stat[13] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[18]~13_combout ;

assign mac_misc_connection_rx_err_stat[14] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[19]~14_combout ;

assign mac_misc_connection_rx_err_stat[15] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[20]~15_combout ;

assign mac_misc_connection_rx_err_stat[16] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[4]~16_combout ;

assign mac_misc_connection_rx_err_stat[17] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_err_stat[22]~17_combout ;

assign mac_misc_connection_rx_frm_type[0] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_ucast~0_combout ;

assign mac_misc_connection_rx_frm_type[1] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_mcast~0_combout ;

assign mac_misc_connection_rx_frm_type[2] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_bcast~0_combout ;

assign mac_misc_connection_rx_frm_type[3] = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|ff_rx_vlan~0_combout ;

assign mac_misc_connection_ff_rx_dsav = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|sav_flag~q ;

assign mac_misc_connection_ff_rx_a_full = \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|afull_flag~q ;

assign mac_misc_connection_ff_rx_a_empty = ~ \eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_RXFF|RX_DATA|aempty_flag~q ;

assign mac_rgmii_connection_rgmii_out[0] = \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[0] ;

assign mac_rgmii_connection_rgmii_out[1] = \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[1] ;

assign mac_rgmii_connection_rgmii_out[2] = \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[2] ;

assign mac_rgmii_connection_rgmii_out[3] = \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out4|altddio_out_component|auto_generated|dataout[3] ;

assign mac_rgmii_connection_tx_control = \eth_tse_0|i_tse_mac|U_RGMII|the_rgmii_out1|altddio_out_component|auto_generated|dataout[0] ;

assign mac_status_connection_eth_mode = \eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|eth_mode~q ;

assign mac_status_connection_ena_10 = \eth_tse_0|i_tse_mac|U_MAC_CONTROL|U_REG|ena_10~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\eth_tse_0|i_tse_mac|U_MAC_TOP|U_MAC|U_TXFF|U_SYNC_2|sync[10].u|std_sync_no_cut|din_s1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFBF7FFFFF7FBFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'h7FFFDFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|AMGP4450_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:1:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:2:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:3:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:4:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:5:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:6:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:7:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:8:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:9:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:10:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:11:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:12:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:13:AMGP4450_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|SQHZ7915:14:AMGP4450_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[10]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[12]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[13]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~1_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal9~0_combout ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[17]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[15]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[16]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|TPOO7242_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|YEAJ1936|JJTX8179[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 .lut_mask = 64'hDEDEDEDEDEDEDEDE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 .lut_mask = 64'hEDDEDEEDDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|BWHK8171_1 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|BWHK8171_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|BWHK8171_2 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|BWHK8171_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|BWHK8171_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|BWHK8171_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|BWHK8171_2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'hDFD5FFFFDFD5FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ZIVV0726~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|FWCA1915[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ZIVV0726~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ZIVV0726 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|ZIVV0726~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|BWHK8171_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ZIVV0726 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|FWCA1915[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|BWHK8171_1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_ZNXJ5711_gen_0:stratixiii_ZNXJ5711_gen_1|ZNXJ5711_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ZIVV0726~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~5_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 .lut_mask = 64'hBFFBFFFFBFFBFFFF;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 .lut_mask = 64'hF9F6F9F6F9F6F9F6;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 .lut_mask = 64'h6996F9F66996F9F6;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~8_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[3]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|VWQM3427|RUGG7005[0]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12 .lut_mask = 64'h7FF7F3777FF7F377;
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113~12_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|VWQM3427|HENC6638~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|FWCA1915[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|FWCA1915[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\altera_internal_jtag~TDIUTAP ),
	.dataf(!\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|sdr (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|sdr .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|sdr .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \nabboc|pzdyqx_impl_inst|sdr .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[11]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[10]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[9]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[8]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[7]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[6]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[5]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[4]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[3]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[2]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[1]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|JJTX8179[0]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|FWCA1915[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VWQM3427|YROJ4113[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|FWCA1915[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|RUWH6717|IHBU8818[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(gnd),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'hCCCCCCCCFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'h66666666FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h55FFAAFF55FFAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h99FF66FF99FF66FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal7~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h69FF96FF69FF96FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 64'h8BFFFFFF8BFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~2_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFAFFFAFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h5F3FFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hAFFAAFFAAFFAAFFA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hBEEBBEEBEBBEEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'hD8FFFFFFD8FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hEFFFFEFFEFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'hFF96FFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hF7FFFFFF37FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

assign \mac_mdio_connection_mdio_in~input_o  = mac_mdio_connection_mdio_in;

endmodule

module IoTOctopus_QSYS_altera_reset_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_32_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_32_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_32_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module IoTOctopus_QSYS_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_IoTOctopus_QSYS_avalon_st_adapter_001 (
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	altera_reset_synchronizer_int_chain_out,
	LessThan0,
	NJQG9082,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	stateLOC_STATE_DATA;
input 	stateLOC_STATE_SHIFT;
input 	altera_reset_synchronizer_int_chain_out;
output 	LessThan0;
input 	NJQG9082;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0 timing_adapter_0(
	.stateLOC_STATE_DATA(stateLOC_STATE_DATA),
	.stateLOC_STATE_SHIFT(stateLOC_STATE_SHIFT),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.LessThan0(LessThan0),
	.NJQG9082(NJQG9082),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0 (
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	altera_reset_synchronizer_int_chain_out,
	LessThan0,
	NJQG9082,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	stateLOC_STATE_DATA;
input 	stateLOC_STATE_SHIFT;
input 	altera_reset_synchronizer_int_chain_out;
output 	LessThan0;
input 	NJQG9082;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[3]~q ;
wire \IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|full~q ;
wire \IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[2]~q ;
wire \IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[1]~q ;
wire \IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[0]~q ;


IoTOctopus_QSYS_IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo_1(
	.stateLOC_STATE_DATA(stateLOC_STATE_DATA),
	.stateLOC_STATE_SHIFT(stateLOC_STATE_SHIFT),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.wr_addr_3(\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[3]~q ),
	.full1(\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|full~q ),
	.wr_addr_2(\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[2]~q ),
	.wr_addr_1(\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[1]~q ),
	.wr_addr_0(\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[0]~q ),
	.NJQG9082(NJQG9082),
	.clk(clk_32_clk));

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[3]~q ),
	.datab(!\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|full~q ),
	.datac(!\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[2]~q ),
	.datad(!\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[1]~q ),
	.datae(!\IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo|wr_addr[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(LessThan0),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_IoTOctopus_QSYS_avalon_st_adapter_001_timing_adapter_0_fifo (
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	reset_n,
	wr_addr_3,
	full1,
	wr_addr_2,
	wr_addr_1,
	wr_addr_0,
	NJQG9082,
	clk)/* synthesis synthesis_greybox=1 */;
input 	stateLOC_STATE_DATA;
input 	stateLOC_STATE_SHIFT;
input 	reset_n;
output 	wr_addr_3;
output 	full1;
output 	wr_addr_2;
output 	wr_addr_1;
output 	wr_addr_0;
input 	NJQG9082;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~0_combout ;
wire \always1~0_combout ;
wire \full~0_combout ;
wire \full~1_combout ;
wire \Add0~1_combout ;
wire \Add0~2_combout ;
wire \wr_addr[0]~0_combout ;


dffeas \wr_addr[3] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(wr_addr_3),
	.prn(vcc));
defparam \wr_addr[3] .is_wysiwyg = "true";
defparam \wr_addr[3] .power_up = "low";

dffeas full(
	.clk(clk),
	.d(\full~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full1),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

dffeas \wr_addr[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(wr_addr_2),
	.prn(vcc));
defparam \wr_addr[2] .is_wysiwyg = "true";
defparam \wr_addr[2] .power_up = "low";

dffeas \wr_addr[1] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(wr_addr_1),
	.prn(vcc));
defparam \wr_addr[1] .is_wysiwyg = "true";
defparam \wr_addr[1] .power_up = "low";

dffeas \wr_addr[0] (
	.clk(clk),
	.d(\wr_addr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(wr_addr_0),
	.prn(vcc));
defparam \wr_addr[0] .is_wysiwyg = "true";
defparam \wr_addr[0] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!wr_addr_3),
	.datab(!wr_addr_2),
	.datac(!wr_addr_1),
	.datad(!wr_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6996699669966996;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!stateLOC_STATE_SHIFT),
	.datab(!stateLOC_STATE_DATA),
	.datac(!NJQG9082),
	.datad(!full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \full~0 (
	.dataa(!wr_addr_3),
	.datab(!wr_addr_2),
	.datac(!wr_addr_1),
	.datad(!wr_addr_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \full~0 .extended_lut = "off";
defparam \full~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \full~0 .shared_arith = "off";

cyclonev_lcell_comb \full~1 (
	.dataa(!stateLOC_STATE_SHIFT),
	.datab(!stateLOC_STATE_DATA),
	.datac(!NJQG9082),
	.datad(!full1),
	.datae(!\full~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \full~1 .extended_lut = "off";
defparam \full~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \full~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!wr_addr_2),
	.datab(!wr_addr_1),
	.datac(!wr_addr_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h9696969696969696;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!wr_addr_1),
	.datab(!wr_addr_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h6666666666666666;
defparam \Add0~2 .shared_arith = "off";

cyclonev_lcell_comb \wr_addr[0]~0 (
	.dataa(!wr_addr_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wr_addr[0]~0 .extended_lut = "off";
defparam \wr_addr[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \wr_addr[0]~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_IoTOctopus_QSYS_eth_tse_0 (
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_01,
	mdio_clk,
	mdio_out,
	command_config_21,
	septy_flag,
	tx_ff_uflow,
	afull_flag,
	aempty_flag,
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	ff_rx_err_stat_5,
	ff_rx_err_stat_6,
	ff_rx_err_stat_7,
	ff_rx_err_stat_8,
	ff_rx_err_stat_9,
	ff_rx_err_stat_10,
	ff_rx_err_stat_11,
	ff_rx_err_stat_12,
	ff_rx_err_stat_13,
	ff_rx_err_stat_14,
	ff_rx_err_stat_15,
	ff_rx_err_stat_16,
	ff_rx_err_stat_17,
	ff_rx_err_stat_18,
	ff_rx_err_stat_19,
	ff_rx_err_stat_20,
	ff_rx_err_stat_4,
	ff_rx_err_stat_22,
	ff_rx_ucast,
	ff_rx_mcast,
	ff_rx_bcast,
	ff_rx_vlan,
	sav_flag,
	afull_flag1,
	aempty_flag1,
	eth_mode,
	ena_10,
	altera_reset_synchronizer_int_chain_out,
	LessThan0,
	din_s1,
	GND_port,
	NJQG9082,
	clk_32_clk,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk,
	mac_status_connection_set_1000,
	mac_status_connection_set_10,
	mac_misc_connection_ff_tx_crc_fwd,
	mac_rgmii_connection_rgmii_in_3,
	mac_rgmii_connection_rgmii_in_2,
	mac_rgmii_connection_rgmii_in_1,
	mac_rgmii_connection_rgmii_in_0,
	mac_rgmii_connection_rx_control,
	mac_misc_connection_magic_sleep_n)/* synthesis synthesis_greybox=1 */;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_01;
output 	mdio_clk;
output 	mdio_out;
output 	command_config_21;
output 	septy_flag;
output 	tx_ff_uflow;
output 	afull_flag;
output 	aempty_flag;
output 	stateLOC_STATE_DATA;
output 	stateLOC_STATE_SHIFT;
output 	ff_rx_err_stat_5;
output 	ff_rx_err_stat_6;
output 	ff_rx_err_stat_7;
output 	ff_rx_err_stat_8;
output 	ff_rx_err_stat_9;
output 	ff_rx_err_stat_10;
output 	ff_rx_err_stat_11;
output 	ff_rx_err_stat_12;
output 	ff_rx_err_stat_13;
output 	ff_rx_err_stat_14;
output 	ff_rx_err_stat_15;
output 	ff_rx_err_stat_16;
output 	ff_rx_err_stat_17;
output 	ff_rx_err_stat_18;
output 	ff_rx_err_stat_19;
output 	ff_rx_err_stat_20;
output 	ff_rx_err_stat_4;
output 	ff_rx_err_stat_22;
output 	ff_rx_ucast;
output 	ff_rx_mcast;
output 	ff_rx_bcast;
output 	ff_rx_vlan;
output 	sav_flag;
output 	afull_flag1;
output 	aempty_flag1;
output 	eth_mode;
output 	ena_10;
input 	altera_reset_synchronizer_int_chain_out;
input 	LessThan0;
output 	din_s1;
input 	GND_port;
input 	NJQG9082;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;
input 	mac_status_connection_set_1000;
input 	mac_status_connection_set_10;
input 	mac_misc_connection_ff_tx_crc_fwd;
input 	mac_rgmii_connection_rgmii_in_3;
input 	mac_rgmii_connection_rgmii_in_2;
input 	mac_rgmii_connection_rgmii_in_1;
input 	mac_rgmii_connection_rgmii_in_0;
input 	mac_rgmii_connection_rx_control;
input 	mac_misc_connection_magic_sleep_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_mac i_tse_mac(
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_01(dataout_01),
	.mdio_clk(mdio_clk),
	.mdio_out(mdio_out),
	.command_config_21(command_config_21),
	.septy_flag(septy_flag),
	.tx_ff_uflow(tx_ff_uflow),
	.afull_flag(afull_flag),
	.aempty_flag(aempty_flag),
	.stateLOC_STATE_DATA(stateLOC_STATE_DATA),
	.stateLOC_STATE_SHIFT(stateLOC_STATE_SHIFT),
	.ff_rx_err_stat_5(ff_rx_err_stat_5),
	.ff_rx_err_stat_6(ff_rx_err_stat_6),
	.ff_rx_err_stat_7(ff_rx_err_stat_7),
	.ff_rx_err_stat_8(ff_rx_err_stat_8),
	.ff_rx_err_stat_9(ff_rx_err_stat_9),
	.ff_rx_err_stat_10(ff_rx_err_stat_10),
	.ff_rx_err_stat_11(ff_rx_err_stat_11),
	.ff_rx_err_stat_12(ff_rx_err_stat_12),
	.ff_rx_err_stat_13(ff_rx_err_stat_13),
	.ff_rx_err_stat_14(ff_rx_err_stat_14),
	.ff_rx_err_stat_15(ff_rx_err_stat_15),
	.ff_rx_err_stat_16(ff_rx_err_stat_16),
	.ff_rx_err_stat_17(ff_rx_err_stat_17),
	.ff_rx_err_stat_18(ff_rx_err_stat_18),
	.ff_rx_err_stat_19(ff_rx_err_stat_19),
	.ff_rx_err_stat_20(ff_rx_err_stat_20),
	.ff_rx_err_stat_4(ff_rx_err_stat_4),
	.ff_rx_err_stat_22(ff_rx_err_stat_22),
	.rx_frm_type({ff_rx_vlan,ff_rx_bcast,ff_rx_mcast,ff_rx_ucast}),
	.sav_flag(sav_flag),
	.afull_flag1(afull_flag1),
	.aempty_flag1(aempty_flag1),
	.eth_mode(eth_mode),
	.ena_10(ena_10),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.LessThan0(LessThan0),
	.din_s1(din_s1),
	.GND_port(GND_port),
	.NJQG9082(NJQG9082),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk),
	.mac_status_connection_set_1000(mac_status_connection_set_1000),
	.mac_status_connection_set_10(mac_status_connection_set_10),
	.mac_misc_connection_ff_tx_crc_fwd(mac_misc_connection_ff_tx_crc_fwd),
	.mac_rgmii_connection_rgmii_in_3(mac_rgmii_connection_rgmii_in_3),
	.mac_rgmii_connection_rgmii_in_2(mac_rgmii_connection_rgmii_in_2),
	.mac_rgmii_connection_rgmii_in_1(mac_rgmii_connection_rgmii_in_1),
	.mac_rgmii_connection_rgmii_in_0(mac_rgmii_connection_rgmii_in_0),
	.mac_rgmii_connection_rx_control(mac_rgmii_connection_rx_control),
	.mac_misc_connection_magic_sleep_n(mac_misc_connection_magic_sleep_n));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_mac (
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_01,
	mdio_clk,
	mdio_out,
	command_config_21,
	septy_flag,
	tx_ff_uflow,
	afull_flag,
	aempty_flag,
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	ff_rx_err_stat_5,
	ff_rx_err_stat_6,
	ff_rx_err_stat_7,
	ff_rx_err_stat_8,
	ff_rx_err_stat_9,
	ff_rx_err_stat_10,
	ff_rx_err_stat_11,
	ff_rx_err_stat_12,
	ff_rx_err_stat_13,
	ff_rx_err_stat_14,
	ff_rx_err_stat_15,
	ff_rx_err_stat_16,
	ff_rx_err_stat_17,
	ff_rx_err_stat_18,
	ff_rx_err_stat_19,
	ff_rx_err_stat_20,
	ff_rx_err_stat_4,
	ff_rx_err_stat_22,
	rx_frm_type,
	sav_flag,
	afull_flag1,
	aempty_flag1,
	eth_mode,
	ena_10,
	altera_reset_synchronizer_int_chain_out,
	LessThan0,
	din_s1,
	GND_port,
	NJQG9082,
	clk_32_clk,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk,
	mac_status_connection_set_1000,
	mac_status_connection_set_10,
	mac_misc_connection_ff_tx_crc_fwd,
	mac_rgmii_connection_rgmii_in_3,
	mac_rgmii_connection_rgmii_in_2,
	mac_rgmii_connection_rgmii_in_1,
	mac_rgmii_connection_rgmii_in_0,
	mac_rgmii_connection_rx_control,
	mac_misc_connection_magic_sleep_n)/* synthesis synthesis_greybox=1 */;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_01;
output 	mdio_clk;
output 	mdio_out;
output 	command_config_21;
output 	septy_flag;
output 	tx_ff_uflow;
output 	afull_flag;
output 	aempty_flag;
output 	stateLOC_STATE_DATA;
output 	stateLOC_STATE_SHIFT;
output 	ff_rx_err_stat_5;
output 	ff_rx_err_stat_6;
output 	ff_rx_err_stat_7;
output 	ff_rx_err_stat_8;
output 	ff_rx_err_stat_9;
output 	ff_rx_err_stat_10;
output 	ff_rx_err_stat_11;
output 	ff_rx_err_stat_12;
output 	ff_rx_err_stat_13;
output 	ff_rx_err_stat_14;
output 	ff_rx_err_stat_15;
output 	ff_rx_err_stat_16;
output 	ff_rx_err_stat_17;
output 	ff_rx_err_stat_18;
output 	ff_rx_err_stat_19;
output 	ff_rx_err_stat_20;
output 	ff_rx_err_stat_4;
output 	ff_rx_err_stat_22;
output 	[3:0] rx_frm_type;
output 	sav_flag;
output 	afull_flag1;
output 	aempty_flag1;
output 	eth_mode;
output 	ena_10;
input 	altera_reset_synchronizer_int_chain_out;
input 	LessThan0;
output 	din_s1;
input 	GND_port;
input 	NJQG9082;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;
input 	mac_status_connection_set_1000;
input 	mac_status_connection_set_10;
input 	mac_misc_connection_ff_tx_crc_fwd;
input 	mac_rgmii_connection_rgmii_in_3;
input 	mac_rgmii_connection_rgmii_in_2;
input 	mac_rgmii_connection_rgmii_in_1;
input 	mac_rgmii_connection_rgmii_in_0;
input 	mac_rgmii_connection_rx_control;
input 	mac_misc_connection_magic_sleep_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[4]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[0]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[5]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[1]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[6]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[2]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[7]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_d_reg[3]~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_err_reg~q ;
wire \U_MAC_TOP|U_GMIF|gm_tx_en_reg~q ;
wire \reset_sync_4|altera_tse_reset_synchronizer_chain_out~q ;
wire \reset_sync_3|altera_tse_reset_synchronizer_chain_out~q ;
wire \reset_sync_1|altera_tse_reset_synchronizer_chain_out~q ;
wire \reset_sync_2|altera_tse_reset_synchronizer_chain_out~q ;
wire \reset_sync_0|altera_tse_reset_synchronizer_chain_out~q ;
wire \U_MAC_TOP|U_MTX|mii_txd_int[0]~q ;
wire \U_MAC_TOP|U_MTX|mii_txd_int[1]~q ;
wire \U_MAC_TOP|U_MTX|mii_txd_int[2]~q ;
wire \U_MAC_TOP|U_MTX|mii_txd_int[3]~q ;
wire \U_MAC_TOP|U_MTX|mii_txerr_int~q ;
wire \U_MAC_TOP|U_MTX|mii_txdv_int~q ;
wire \U_MAC_TOP|U_MAC|U_MAGIC|magic_detect~q ;
wire \U_MAC_CONTROL|U_REG|ethernet_mode~q ;
wire \U_MAC_CONTROL|U_REG|sleep_ena~q ;
wire \U_RGMII|U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \U_RGMII|rx_dv~q ;
wire \U_RGMII|rgmii_in_4_reg[7]~q ;
wire \U_RGMII|rgmii_in_4_reg[6]~q ;
wire \U_RGMII|rgmii_in_4_reg[5]~q ;
wire \U_RGMII|rgmii_in_4_reg[4]~q ;
wire \U_RGMII|rgmii_in_4_reg[0]~q ;
wire \U_RGMII|rgmii_in_4_reg[3]~q ;
wire \U_RGMII|rgmii_in_4_reg[2]~q ;
wire \U_RGMII|rgmii_in_4_reg[1]~q ;
wire \U_RGMII|m_rx_crs~2_combout ;
wire \U_MAC_TOP|neinyesfmd~55_combout ;
wire \U_RGMII|gm_rx_err~combout ;


IoTOctopus_QSYS_altera_tse_top_w_fifo_10_100_1000 U_MAC_TOP(
	.gm_tx_d_reg_4(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[4]~q ),
	.gm_tx_d_reg_0(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[0]~q ),
	.gm_tx_d_reg_5(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[5]~q ),
	.gm_tx_d_reg_1(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[1]~q ),
	.gm_tx_d_reg_6(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[6]~q ),
	.gm_tx_d_reg_2(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[2]~q ),
	.gm_tx_d_reg_7(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[7]~q ),
	.gm_tx_d_reg_3(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[3]~q ),
	.gm_tx_err_reg(\U_MAC_TOP|U_GMIF|gm_tx_err_reg~q ),
	.gm_tx_en_reg(\U_MAC_TOP|U_GMIF|gm_tx_en_reg~q ),
	.septy_flag(septy_flag),
	.tx_ff_uflow(tx_ff_uflow),
	.afull_flag(afull_flag),
	.aempty_flag(aempty_flag),
	.stateLOC_STATE_DATA(stateLOC_STATE_DATA),
	.stateLOC_STATE_SHIFT(stateLOC_STATE_SHIFT),
	.ff_rx_err_stat_5(ff_rx_err_stat_5),
	.ff_rx_err_stat_6(ff_rx_err_stat_6),
	.ff_rx_err_stat_7(ff_rx_err_stat_7),
	.ff_rx_err_stat_8(ff_rx_err_stat_8),
	.ff_rx_err_stat_9(ff_rx_err_stat_9),
	.ff_rx_err_stat_10(ff_rx_err_stat_10),
	.ff_rx_err_stat_11(ff_rx_err_stat_11),
	.ff_rx_err_stat_12(ff_rx_err_stat_12),
	.ff_rx_err_stat_13(ff_rx_err_stat_13),
	.ff_rx_err_stat_14(ff_rx_err_stat_14),
	.ff_rx_err_stat_15(ff_rx_err_stat_15),
	.ff_rx_err_stat_16(ff_rx_err_stat_16),
	.ff_rx_err_stat_17(ff_rx_err_stat_17),
	.ff_rx_err_stat_18(ff_rx_err_stat_18),
	.ff_rx_err_stat_19(ff_rx_err_stat_19),
	.ff_rx_err_stat_20(ff_rx_err_stat_20),
	.ff_rx_err_stat_4(ff_rx_err_stat_4),
	.ff_rx_err_stat_22(ff_rx_err_stat_22),
	.ff_rx_ucast(rx_frm_type[0]),
	.ff_rx_mcast(rx_frm_type[1]),
	.ff_rx_bcast(rx_frm_type[2]),
	.ff_rx_vlan(rx_frm_type[3]),
	.sav_flag(sav_flag),
	.afull_flag1(afull_flag1),
	.aempty_flag1(aempty_flag1),
	.altera_tse_reset_synchronizer_chain_out(\reset_sync_3|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_tse_reset_synchronizer_chain_out1(\reset_sync_1|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_tse_reset_synchronizer_chain_out2(\reset_sync_2|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_tse_reset_synchronizer_chain_out3(\reset_sync_0|altera_tse_reset_synchronizer_chain_out~q ),
	.mii_txd_int_0(\U_MAC_TOP|U_MTX|mii_txd_int[0]~q ),
	.mii_txd_int_1(\U_MAC_TOP|U_MTX|mii_txd_int[1]~q ),
	.mii_txd_int_2(\U_MAC_TOP|U_MTX|mii_txd_int[2]~q ),
	.mii_txd_int_3(\U_MAC_TOP|U_MTX|mii_txd_int[3]~q ),
	.mii_txerr_int(\U_MAC_TOP|U_MTX|mii_txerr_int~q ),
	.mii_txdv_int(\U_MAC_TOP|U_MTX|mii_txdv_int~q ),
	.LessThan0(LessThan0),
	.magic_detect(\U_MAC_TOP|U_MAC|U_MAGIC|magic_detect~q ),
	.ethernet_mode(\U_MAC_CONTROL|U_REG|ethernet_mode~q ),
	.sleep_ena(\U_MAC_CONTROL|U_REG|sleep_ena~q ),
	.dreg_1(\U_RGMII|U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.rx_dv(\U_RGMII|rx_dv~q ),
	.rgmii_in_4_reg_7(\U_RGMII|rgmii_in_4_reg[7]~q ),
	.rgmii_in_4_reg_6(\U_RGMII|rgmii_in_4_reg[6]~q ),
	.rgmii_in_4_reg_5(\U_RGMII|rgmii_in_4_reg[5]~q ),
	.rgmii_in_4_reg_4(\U_RGMII|rgmii_in_4_reg[4]~q ),
	.rgmii_in_4_reg_0(\U_RGMII|rgmii_in_4_reg[0]~q ),
	.rgmii_in_4_reg_3(\U_RGMII|rgmii_in_4_reg[3]~q ),
	.rgmii_in_4_reg_2(\U_RGMII|rgmii_in_4_reg[2]~q ),
	.rgmii_in_4_reg_1(\U_RGMII|rgmii_in_4_reg[1]~q ),
	.m_rx_crs(\U_RGMII|m_rx_crs~2_combout ),
	.neinyesfmd(\U_MAC_TOP|neinyesfmd~55_combout ),
	.gm_rx_err(\U_RGMII|gm_rx_err~combout ),
	.din_s1(din_s1),
	.GND_port(GND_port),
	.NJQG9082(NJQG9082),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk),
	.mac_misc_connection_ff_tx_crc_fwd(mac_misc_connection_ff_tx_crc_fwd));

IoTOctopus_QSYS_altera_tse_rgmii_module U_RGMII(
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.dataout_01(dataout_01),
	.gm_tx_d_reg_4(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[4]~q ),
	.gm_tx_d_reg_0(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[0]~q ),
	.gm_tx_d_reg_5(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[5]~q ),
	.gm_tx_d_reg_1(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[1]~q ),
	.gm_tx_d_reg_6(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[6]~q ),
	.gm_tx_d_reg_2(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[2]~q ),
	.gm_tx_d_reg_7(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[7]~q ),
	.gm_tx_d_reg_3(\U_MAC_TOP|U_GMIF|gm_tx_d_reg[3]~q ),
	.gm_tx_err_reg(\U_MAC_TOP|U_GMIF|gm_tx_err_reg~q ),
	.gm_tx_en_reg(\U_MAC_TOP|U_GMIF|gm_tx_en_reg~q ),
	.eth_mode(eth_mode),
	.altera_tse_reset_synchronizer_chain_out(\reset_sync_1|altera_tse_reset_synchronizer_chain_out~q ),
	.reset_rx_clk(\reset_sync_0|altera_tse_reset_synchronizer_chain_out~q ),
	.mii_txd_int_0(\U_MAC_TOP|U_MTX|mii_txd_int[0]~q ),
	.mii_txd_int_1(\U_MAC_TOP|U_MTX|mii_txd_int[1]~q ),
	.mii_txd_int_2(\U_MAC_TOP|U_MTX|mii_txd_int[2]~q ),
	.mii_txd_int_3(\U_MAC_TOP|U_MTX|mii_txd_int[3]~q ),
	.mii_txerr_int(\U_MAC_TOP|U_MTX|mii_txerr_int~q ),
	.mii_txdv_int(\U_MAC_TOP|U_MTX|mii_txdv_int~q ),
	.dreg_1(\U_RGMII|U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.rx_dv1(\U_RGMII|rx_dv~q ),
	.rgmii_in_4_reg_7(\U_RGMII|rgmii_in_4_reg[7]~q ),
	.rgmii_in_4_reg_6(\U_RGMII|rgmii_in_4_reg[6]~q ),
	.rgmii_in_4_reg_5(\U_RGMII|rgmii_in_4_reg[5]~q ),
	.rgmii_in_4_reg_4(\U_RGMII|rgmii_in_4_reg[4]~q ),
	.rgmii_in_4_reg_0(\U_RGMII|rgmii_in_4_reg[0]~q ),
	.rgmii_in_4_reg_3(\U_RGMII|rgmii_in_4_reg[3]~q ),
	.rgmii_in_4_reg_2(\U_RGMII|rgmii_in_4_reg[2]~q ),
	.rgmii_in_4_reg_1(\U_RGMII|rgmii_in_4_reg[1]~q ),
	.m_rx_crs(\U_RGMII|m_rx_crs~2_combout ),
	.m_tx_en(\U_MAC_TOP|neinyesfmd~55_combout ),
	.gm_rx_err1(\U_RGMII|gm_rx_err~combout ),
	.NJQG9082(NJQG9082),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk),
	.mac_rgmii_connection_rgmii_in_3(mac_rgmii_connection_rgmii_in_3),
	.mac_rgmii_connection_rgmii_in_2(mac_rgmii_connection_rgmii_in_2),
	.mac_rgmii_connection_rgmii_in_1(mac_rgmii_connection_rgmii_in_1),
	.mac_rgmii_connection_rgmii_in_0(mac_rgmii_connection_rgmii_in_0),
	.mac_rgmii_connection_rx_control(mac_rgmii_connection_rx_control));

IoTOctopus_QSYS_altera_tse_top_mdio U_MDIO(
	.mdio_clk(mdio_clk),
	.mdio_out1(mdio_out),
	.altera_tse_reset_synchronizer_chain_out(\reset_sync_4|altera_tse_reset_synchronizer_chain_out~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_mac_control U_MAC_CONTROL(
	.command_config_21(command_config_21),
	.eth_mode(eth_mode),
	.ena_10(ena_10),
	.altera_tse_reset_synchronizer_chain_out(\reset_sync_4|altera_tse_reset_synchronizer_chain_out~q ),
	.magic_detect(\U_MAC_TOP|U_MAC|U_MAGIC|magic_detect~q ),
	.ethernet_mode(\U_MAC_CONTROL|U_REG|ethernet_mode~q ),
	.sleep_ena(\U_MAC_CONTROL|U_REG|sleep_ena~q ),
	.clk_32_clk(clk_32_clk),
	.mac_status_connection_set_1000(mac_status_connection_set_1000),
	.mac_status_connection_set_10(mac_status_connection_set_10),
	.mac_misc_connection_magic_sleep_n(mac_misc_connection_magic_sleep_n));

IoTOctopus_QSYS_altera_tse_reset_synchronizer_4 reset_sync_4(
	.altera_tse_reset_synchronizer_chain_out1(\reset_sync_4|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_reset_synchronizer_3 reset_sync_3(
	.altera_tse_reset_synchronizer_chain_out1(\reset_sync_3|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_reset_synchronizer_2 reset_sync_2(
	.altera_tse_reset_synchronizer_chain_out1(\reset_sync_2|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_reset_synchronizer_1 reset_sync_1(
	.altera_tse_reset_synchronizer_chain_out1(\reset_sync_1|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_reset_synchronizer reset_sync_0(
	.altera_tse_reset_synchronizer_chain_out1(\reset_sync_0|altera_tse_reset_synchronizer_chain_out~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_tse_mac_control (
	command_config_21,
	eth_mode,
	ena_10,
	altera_tse_reset_synchronizer_chain_out,
	magic_detect,
	ethernet_mode,
	sleep_ena,
	clk_32_clk,
	mac_status_connection_set_1000,
	mac_status_connection_set_10,
	mac_misc_connection_magic_sleep_n)/* synthesis synthesis_greybox=1 */;
output 	command_config_21;
output 	eth_mode;
output 	ena_10;
input 	altera_tse_reset_synchronizer_chain_out;
input 	magic_detect;
output 	ethernet_mode;
output 	sleep_ena;
input 	clk_32_clk;
input 	mac_status_connection_set_1000;
input 	mac_status_connection_set_10;
input 	mac_misc_connection_magic_sleep_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_tse_register_map U_REG(
	.command_config_21(command_config_21),
	.eth_mode1(eth_mode),
	.ena_101(ena_10),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.magic_detect(magic_detect),
	.ethernet_mode1(ethernet_mode),
	.sleep_ena1(sleep_ena),
	.clk_32_clk(clk_32_clk),
	.mac_status_connection_set_1000(mac_status_connection_set_1000),
	.mac_status_connection_set_10(mac_status_connection_set_10),
	.mac_misc_connection_magic_sleep_n(mac_misc_connection_magic_sleep_n));

endmodule

module IoTOctopus_QSYS_altera_tse_register_map (
	command_config_21,
	eth_mode1,
	ena_101,
	altera_tse_reset_synchronizer_chain_out,
	magic_detect,
	ethernet_mode1,
	sleep_ena1,
	clk_32_clk,
	mac_status_connection_set_1000,
	mac_status_connection_set_10,
	mac_misc_connection_magic_sleep_n)/* synthesis synthesis_greybox=1 */;
output 	command_config_21;
output 	eth_mode1;
output 	ena_101;
input 	altera_tse_reset_synchronizer_chain_out;
input 	magic_detect;
output 	ethernet_mode1;
output 	sleep_ena1;
input 	clk_32_clk;
input 	mac_status_connection_set_1000;
input 	mac_status_connection_set_10;
input 	mac_misc_connection_magic_sleep_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_MAGIC_DETECT|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \sleep_ena~0_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_2 U_MAGIC_DETECT(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_MAGIC_DETECT|std_sync_no_cut|dreg[1]~q ),
	.magic_detect(magic_detect),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_3 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk),
	.mac_misc_connection_magic_sleep_n(mac_misc_connection_magic_sleep_n));

dffeas \command_config[21] (
	.clk(clk_32_clk),
	.d(\U_MAGIC_DETECT|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(command_config_21),
	.prn(vcc));
defparam \command_config[21] .is_wysiwyg = "true";
defparam \command_config[21] .power_up = "low";

dffeas eth_mode(
	.clk(clk_32_clk),
	.d(mac_status_connection_set_1000),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(eth_mode1),
	.prn(vcc));
defparam eth_mode.is_wysiwyg = "true";
defparam eth_mode.power_up = "low";

dffeas ena_10(
	.clk(clk_32_clk),
	.d(mac_status_connection_set_10),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ena_101),
	.prn(vcc));
defparam ena_10.is_wysiwyg = "true";
defparam ena_10.power_up = "low";

dffeas ethernet_mode(
	.clk(clk_32_clk),
	.d(mac_status_connection_set_1000),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ethernet_mode1),
	.prn(vcc));
defparam ethernet_mode.is_wysiwyg = "true";
defparam ethernet_mode.power_up = "low";

dffeas sleep_ena(
	.clk(clk_32_clk),
	.d(\sleep_ena~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sleep_ena1),
	.prn(vcc));
defparam sleep_ena.is_wysiwyg = "true";
defparam sleep_ena.power_up = "low";

cyclonev_lcell_comb \sleep_ena~0 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sleep_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sleep_ena~0 .extended_lut = "off";
defparam \sleep_ena~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \sleep_ena~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_2 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	magic_detect,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	magic_detect;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_2 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(magic_detect),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_2 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_3 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk,
	mac_misc_connection_magic_sleep_n)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;
input 	mac_misc_connection_magic_sleep_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_5 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk),
	.din(mac_misc_connection_magic_sleep_n));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_5 (
	reset_n,
	dreg_1,
	clk,
	din)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;
input 	din;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_reset_synchronizer (
	altera_tse_reset_synchronizer_chain_out1,
	altera_reset_synchronizer_int_chain_out,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_tse_reset_synchronizer_chain[1]~q ;
wire \altera_tse_reset_synchronizer_chain[0]~q ;


dffeas altera_tse_reset_synchronizer_chain_out(
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_tse_reset_synchronizer_chain_out1),
	.prn(vcc));
defparam altera_tse_reset_synchronizer_chain_out.is_wysiwyg = "true";
defparam altera_tse_reset_synchronizer_chain_out.power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[1]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[1] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[1] .power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[0] (
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[0]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[0] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_reset_synchronizer_1 (
	altera_tse_reset_synchronizer_chain_out1,
	altera_reset_synchronizer_int_chain_out,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_tse_reset_synchronizer_chain[1]~q ;
wire \altera_tse_reset_synchronizer_chain[0]~q ;


dffeas altera_tse_reset_synchronizer_chain_out(
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_tse_reset_synchronizer_chain_out1),
	.prn(vcc));
defparam altera_tse_reset_synchronizer_chain_out.is_wysiwyg = "true";
defparam altera_tse_reset_synchronizer_chain_out.power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[1]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[1] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[1] .power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[0] (
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[0]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[0] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_reset_synchronizer_2 (
	altera_tse_reset_synchronizer_chain_out1,
	altera_reset_synchronizer_int_chain_out,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_tse_reset_synchronizer_chain[1]~q ;
wire \altera_tse_reset_synchronizer_chain[0]~q ;


dffeas altera_tse_reset_synchronizer_chain_out(
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_tse_reset_synchronizer_chain_out1),
	.prn(vcc));
defparam altera_tse_reset_synchronizer_chain_out.is_wysiwyg = "true";
defparam altera_tse_reset_synchronizer_chain_out.power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[1]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[1] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[1] .power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[0] (
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[0]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[0] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_reset_synchronizer_3 (
	altera_tse_reset_synchronizer_chain_out1,
	altera_reset_synchronizer_int_chain_out,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_tse_reset_synchronizer_chain[1]~q ;
wire \altera_tse_reset_synchronizer_chain[0]~q ;


dffeas altera_tse_reset_synchronizer_chain_out(
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_tse_reset_synchronizer_chain_out1),
	.prn(vcc));
defparam altera_tse_reset_synchronizer_chain_out.is_wysiwyg = "true";
defparam altera_tse_reset_synchronizer_chain_out.power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[1]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[1] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[1] .power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[0] (
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[0]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[0] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_reset_synchronizer_4 (
	altera_tse_reset_synchronizer_chain_out1,
	altera_reset_synchronizer_int_chain_out,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_tse_reset_synchronizer_chain[1]~q ;
wire \altera_tse_reset_synchronizer_chain[0]~q ;


dffeas altera_tse_reset_synchronizer_chain_out(
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_tse_reset_synchronizer_chain_out1),
	.prn(vcc));
defparam altera_tse_reset_synchronizer_chain_out.is_wysiwyg = "true";
defparam altera_tse_reset_synchronizer_chain_out.power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[1]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[1] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[1] .power_up = "low";

dffeas \altera_tse_reset_synchronizer_chain[0] (
	.clk(clk),
	.d(\altera_tse_reset_synchronizer_chain[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_tse_reset_synchronizer_chain[0]~q ),
	.prn(vcc));
defparam \altera_tse_reset_synchronizer_chain[0] .is_wysiwyg = "true";
defparam \altera_tse_reset_synchronizer_chain[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_rgmii_module (
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	dataout_01,
	gm_tx_d_reg_4,
	gm_tx_d_reg_0,
	gm_tx_d_reg_5,
	gm_tx_d_reg_1,
	gm_tx_d_reg_6,
	gm_tx_d_reg_2,
	gm_tx_d_reg_7,
	gm_tx_d_reg_3,
	gm_tx_err_reg,
	gm_tx_en_reg,
	eth_mode,
	altera_tse_reset_synchronizer_chain_out,
	reset_rx_clk,
	mii_txd_int_0,
	mii_txd_int_1,
	mii_txd_int_2,
	mii_txd_int_3,
	mii_txerr_int,
	mii_txdv_int,
	dreg_1,
	rx_dv1,
	rgmii_in_4_reg_7,
	rgmii_in_4_reg_6,
	rgmii_in_4_reg_5,
	rgmii_in_4_reg_4,
	rgmii_in_4_reg_0,
	rgmii_in_4_reg_3,
	rgmii_in_4_reg_2,
	rgmii_in_4_reg_1,
	m_rx_crs,
	m_tx_en,
	gm_rx_err1,
	NJQG9082,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk,
	mac_rgmii_connection_rgmii_in_3,
	mac_rgmii_connection_rgmii_in_2,
	mac_rgmii_connection_rgmii_in_1,
	mac_rgmii_connection_rgmii_in_0,
	mac_rgmii_connection_rx_control)/* synthesis synthesis_greybox=1 */;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
output 	dataout_01;
input 	gm_tx_d_reg_4;
input 	gm_tx_d_reg_0;
input 	gm_tx_d_reg_5;
input 	gm_tx_d_reg_1;
input 	gm_tx_d_reg_6;
input 	gm_tx_d_reg_2;
input 	gm_tx_d_reg_7;
input 	gm_tx_d_reg_3;
input 	gm_tx_err_reg;
input 	gm_tx_en_reg;
input 	eth_mode;
input 	altera_tse_reset_synchronizer_chain_out;
input 	reset_rx_clk;
input 	mii_txd_int_0;
input 	mii_txd_int_1;
input 	mii_txd_int_2;
input 	mii_txd_int_3;
input 	mii_txerr_int;
input 	mii_txdv_int;
output 	dreg_1;
output 	rx_dv1;
output 	rgmii_in_4_reg_7;
output 	rgmii_in_4_reg_6;
output 	rgmii_in_4_reg_5;
output 	rgmii_in_4_reg_4;
output 	rgmii_in_4_reg_0;
output 	rgmii_in_4_reg_3;
output 	rgmii_in_4_reg_2;
output 	rgmii_in_4_reg_1;
output 	m_rx_crs;
input 	m_tx_en;
output 	gm_rx_err1;
input 	NJQG9082;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;
input 	mac_rgmii_connection_rgmii_in_3;
input 	mac_rgmii_connection_rgmii_in_2;
input 	mac_rgmii_connection_rgmii_in_1;
input 	mac_rgmii_connection_rgmii_in_0;
input 	mac_rgmii_connection_rx_control;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[3] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[3] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[2] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[2] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[1] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[1] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[0] ;
wire \the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[0] ;
wire \the_rgmii_in1|altddio_in_component|auto_generated|dataout_l[0] ;
wire \the_rgmii_in1|altddio_in_component|auto_generated|dataout_h[0] ;
wire \U_SYNC_2|std_sync_no_cut|dreg[1]~q ;
wire \rgmii_out_4_wire[4]~0_combout ;
wire \rgmii_out_4_wire[0]~1_combout ;
wire \rgmii_out_4_wire[5]~2_combout ;
wire \rgmii_out_4_wire[1]~3_combout ;
wire \rgmii_out_4_wire[6]~4_combout ;
wire \rgmii_out_4_wire[2]~5_combout ;
wire \rgmii_out_4_wire[7]~6_combout ;
wire \rgmii_out_4_wire[3]~7_combout ;
wire \rgmii_out_1_wire_inp2~0_combout ;
wire \rgmii_out_1_wire_inp1~0_combout ;
wire \m_tx_en_reg4~q ;
wire \m_rx_col_reg~0_combout ;
wire \m_tx_en_reg3~q ;
wire \m_tx_en_reg2~q ;
wire \m_tx_en_reg1~q ;
wire \rgmii_in_1_temp_reg[1]~q ;
wire \rgmii_in_4_temp_reg[4]~q ;
wire \rgmii_in_4_temp_reg[7]~q ;
wire \rgmii_in_4_temp_reg[6]~q ;
wire \rgmii_in_4_temp_reg[5]~q ;
wire \m_rx_crs~0_combout ;
wire \rx_err~q ;
wire \m_rx_crs~1_combout ;


IoTOctopus_QSYS_altera_tse_rgmii_out1 the_rgmii_out1(
	.dataout_0(dataout_01),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.rgmii_out_1_wire_inp2(\rgmii_out_1_wire_inp2~0_combout ),
	.rgmii_out_1_wire_inp1(\rgmii_out_1_wire_inp1~0_combout ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_rgmii_out4 the_rgmii_out4(
	.dataout_0(dataout_0),
	.dataout_1(dataout_1),
	.dataout_2(dataout_2),
	.dataout_3(dataout_3),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.rgmii_out_4_wire_4(\rgmii_out_4_wire[4]~0_combout ),
	.rgmii_out_4_wire_0(\rgmii_out_4_wire[0]~1_combout ),
	.rgmii_out_4_wire_5(\rgmii_out_4_wire[5]~2_combout ),
	.rgmii_out_4_wire_1(\rgmii_out_4_wire[1]~3_combout ),
	.rgmii_out_4_wire_6(\rgmii_out_4_wire[6]~4_combout ),
	.rgmii_out_4_wire_2(\rgmii_out_4_wire[2]~5_combout ),
	.rgmii_out_4_wire_7(\rgmii_out_4_wire[7]~6_combout ),
	.rgmii_out_4_wire_3(\rgmii_out_4_wire[3]~7_combout ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_15 U_SYNC_2(
	.eth_mode(eth_mode),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_14 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.m_rx_col_reg(\m_rx_col_reg~0_combout ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_rgmii_in1 the_rgmii_in1(
	.dataout_l_0(\the_rgmii_in1|altddio_in_component|auto_generated|dataout_l[0] ),
	.dataout_h_0(\the_rgmii_in1|altddio_in_component|auto_generated|dataout_h[0] ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk),
	.mac_rgmii_connection_rx_control(mac_rgmii_connection_rx_control));

IoTOctopus_QSYS_altera_tse_rgmii_in4 the_rgmii_in4(
	.dataout_l_3(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[3] ),
	.dataout_h_3(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[3] ),
	.dataout_l_2(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[2] ),
	.dataout_h_2(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[2] ),
	.dataout_l_1(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[1] ),
	.dataout_h_1(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[1] ),
	.dataout_l_0(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[0] ),
	.dataout_h_0(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[0] ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk),
	.mac_rgmii_connection_rgmii_in_3(mac_rgmii_connection_rgmii_in_3),
	.mac_rgmii_connection_rgmii_in_2(mac_rgmii_connection_rgmii_in_2),
	.mac_rgmii_connection_rgmii_in_1(mac_rgmii_connection_rgmii_in_1),
	.mac_rgmii_connection_rgmii_in_0(mac_rgmii_connection_rgmii_in_0));

cyclonev_lcell_comb \rgmii_out_4_wire[4]~0 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!gm_tx_d_reg_4),
	.datad(!mii_txd_int_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[4]~0 .extended_lut = "off";
defparam \rgmii_out_4_wire[4]~0 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[0]~1 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!mii_txd_int_0),
	.datad(!gm_tx_d_reg_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[0]~1 .extended_lut = "off";
defparam \rgmii_out_4_wire[0]~1 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[5]~2 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!gm_tx_d_reg_5),
	.datad(!mii_txd_int_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[5]~2 .extended_lut = "off";
defparam \rgmii_out_4_wire[5]~2 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[1]~3 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!mii_txd_int_1),
	.datad(!gm_tx_d_reg_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[1]~3 .extended_lut = "off";
defparam \rgmii_out_4_wire[1]~3 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[6]~4 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!gm_tx_d_reg_6),
	.datad(!mii_txd_int_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[6]~4 .extended_lut = "off";
defparam \rgmii_out_4_wire[6]~4 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[2]~5 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!mii_txd_int_2),
	.datad(!gm_tx_d_reg_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[2]~5 .extended_lut = "off";
defparam \rgmii_out_4_wire[2]~5 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[7]~6 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!gm_tx_d_reg_7),
	.datad(!mii_txd_int_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[7]~6 .extended_lut = "off";
defparam \rgmii_out_4_wire[7]~6 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[7]~6 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_4_wire[3]~7 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!mii_txd_int_3),
	.datad(!gm_tx_d_reg_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_4_wire[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_4_wire[3]~7 .extended_lut = "off";
defparam \rgmii_out_4_wire[3]~7 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_4_wire[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_1_wire_inp2~0 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!gm_tx_err_reg),
	.datad(!gm_tx_en_reg),
	.datae(!mii_txerr_int),
	.dataf(!mii_txdv_int),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_1_wire_inp2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_1_wire_inp2~0 .extended_lut = "off";
defparam \rgmii_out_1_wire_inp2~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \rgmii_out_1_wire_inp2~0 .shared_arith = "off";

cyclonev_lcell_comb \rgmii_out_1_wire_inp1~0 (
	.dataa(!NJQG9082),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(!gm_tx_en_reg),
	.datad(!mii_txdv_int),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rgmii_out_1_wire_inp1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rgmii_out_1_wire_inp1~0 .extended_lut = "off";
defparam \rgmii_out_1_wire_inp1~0 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \rgmii_out_1_wire_inp1~0 .shared_arith = "off";

dffeas m_tx_en_reg4(
	.clk(mac_tx_clock_connection_clk),
	.d(\m_tx_en_reg3~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_tx_en_reg4~q ),
	.prn(vcc));
defparam m_tx_en_reg4.is_wysiwyg = "true";
defparam m_tx_en_reg4.power_up = "low";

cyclonev_lcell_comb \m_rx_col_reg~0 (
	.dataa(!rx_dv1),
	.datab(!\m_rx_crs~0_combout ),
	.datac(!\m_rx_crs~1_combout ),
	.datad(!\m_tx_en_reg4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_rx_col_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_rx_col_reg~0 .extended_lut = "off";
defparam \m_rx_col_reg~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \m_rx_col_reg~0 .shared_arith = "off";

dffeas m_tx_en_reg3(
	.clk(mac_tx_clock_connection_clk),
	.d(\m_tx_en_reg2~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_tx_en_reg3~q ),
	.prn(vcc));
defparam m_tx_en_reg3.is_wysiwyg = "true";
defparam m_tx_en_reg3.power_up = "low";

dffeas m_tx_en_reg2(
	.clk(mac_tx_clock_connection_clk),
	.d(\m_tx_en_reg1~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_tx_en_reg2~q ),
	.prn(vcc));
defparam m_tx_en_reg2.is_wysiwyg = "true";
defparam m_tx_en_reg2.power_up = "low";

dffeas m_tx_en_reg1(
	.clk(mac_tx_clock_connection_clk),
	.d(m_tx_en),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\m_tx_en_reg1~q ),
	.prn(vcc));
defparam m_tx_en_reg1.is_wysiwyg = "true";
defparam m_tx_en_reg1.power_up = "low";

dffeas rx_dv(
	.clk(mac_rx_clock_connection_clk),
	.d(\rgmii_in_1_temp_reg[1]~q ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_dv1),
	.prn(vcc));
defparam rx_dv.is_wysiwyg = "true";
defparam rx_dv.power_up = "low";

dffeas \rgmii_in_4_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[3] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_7),
	.prn(vcc));
defparam \rgmii_in_4_reg[7] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[7] .power_up = "low";

dffeas \rgmii_in_4_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[2] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_6),
	.prn(vcc));
defparam \rgmii_in_4_reg[6] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[6] .power_up = "low";

dffeas \rgmii_in_4_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[1] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_5),
	.prn(vcc));
defparam \rgmii_in_4_reg[5] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[5] .power_up = "low";

dffeas \rgmii_in_4_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_l[0] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_4),
	.prn(vcc));
defparam \rgmii_in_4_reg[4] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[4] .power_up = "low";

dffeas \rgmii_in_4_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rgmii_in_4_temp_reg[4]~q ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_0),
	.prn(vcc));
defparam \rgmii_in_4_reg[0] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[0] .power_up = "low";

dffeas \rgmii_in_4_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rgmii_in_4_temp_reg[7]~q ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_3),
	.prn(vcc));
defparam \rgmii_in_4_reg[3] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[3] .power_up = "low";

dffeas \rgmii_in_4_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rgmii_in_4_temp_reg[6]~q ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_2),
	.prn(vcc));
defparam \rgmii_in_4_reg[2] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[2] .power_up = "low";

dffeas \rgmii_in_4_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rgmii_in_4_temp_reg[5]~q ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rgmii_in_4_reg_1),
	.prn(vcc));
defparam \rgmii_in_4_reg[1] .is_wysiwyg = "true";
defparam \rgmii_in_4_reg[1] .power_up = "low";

cyclonev_lcell_comb \m_rx_crs~2 (
	.dataa(!rx_dv1),
	.datab(!\m_rx_crs~0_combout ),
	.datac(!\m_rx_crs~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m_rx_crs),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_rx_crs~2 .extended_lut = "off";
defparam \m_rx_crs~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \m_rx_crs~2 .shared_arith = "off";

cyclonev_lcell_comb gm_rx_err(
	.dataa(!rx_dv1),
	.datab(!\rx_err~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(gm_rx_err1),
	.sumout(),
	.cout(),
	.shareout());
defparam gm_rx_err.extended_lut = "off";
defparam gm_rx_err.lut_mask = 64'h6666666666666666;
defparam gm_rx_err.shared_arith = "off";

dffeas \rgmii_in_1_temp_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in1|altddio_in_component|auto_generated|dataout_h[0] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rgmii_in_1_temp_reg[1]~q ),
	.prn(vcc));
defparam \rgmii_in_1_temp_reg[1] .is_wysiwyg = "true";
defparam \rgmii_in_1_temp_reg[1] .power_up = "low";

dffeas \rgmii_in_4_temp_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[0] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rgmii_in_4_temp_reg[4]~q ),
	.prn(vcc));
defparam \rgmii_in_4_temp_reg[4] .is_wysiwyg = "true";
defparam \rgmii_in_4_temp_reg[4] .power_up = "low";

dffeas \rgmii_in_4_temp_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[3] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rgmii_in_4_temp_reg[7]~q ),
	.prn(vcc));
defparam \rgmii_in_4_temp_reg[7] .is_wysiwyg = "true";
defparam \rgmii_in_4_temp_reg[7] .power_up = "low";

dffeas \rgmii_in_4_temp_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[2] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rgmii_in_4_temp_reg[6]~q ),
	.prn(vcc));
defparam \rgmii_in_4_temp_reg[6] .is_wysiwyg = "true";
defparam \rgmii_in_4_temp_reg[6] .power_up = "low";

dffeas \rgmii_in_4_temp_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in4|altddio_in_component|auto_generated|dataout_h[1] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rgmii_in_4_temp_reg[5]~q ),
	.prn(vcc));
defparam \rgmii_in_4_temp_reg[5] .is_wysiwyg = "true";
defparam \rgmii_in_4_temp_reg[5] .power_up = "low";

cyclonev_lcell_comb \m_rx_crs~0 (
	.dataa(!rgmii_in_4_reg_7),
	.datab(!rgmii_in_4_reg_6),
	.datac(!rgmii_in_4_reg_5),
	.datad(!rgmii_in_4_reg_4),
	.datae(!rgmii_in_4_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_rx_crs~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_rx_crs~0 .extended_lut = "off";
defparam \m_rx_crs~0 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \m_rx_crs~0 .shared_arith = "off";

dffeas rx_err(
	.clk(mac_rx_clock_connection_clk),
	.d(\the_rgmii_in1|altddio_in_component|auto_generated|dataout_l[0] ),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rx_err~q ),
	.prn(vcc));
defparam rx_err.is_wysiwyg = "true";
defparam rx_err.power_up = "low";

cyclonev_lcell_comb \m_rx_crs~1 (
	.dataa(!rgmii_in_4_reg_3),
	.datab(!rgmii_in_4_reg_2),
	.datac(!rgmii_in_4_reg_1),
	.datad(!\rx_err~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\m_rx_crs~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \m_rx_crs~1 .extended_lut = "off";
defparam \m_rx_crs~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \m_rx_crs~1 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_14 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	m_rx_col_reg,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	m_rx_col_reg;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_14 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(m_rx_col_reg),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_14 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_15 (
	eth_mode,
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	eth_mode;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_15 std_sync_no_cut(
	.din(eth_mode),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_15 (
	din,
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_rgmii_in1 (
	dataout_l_0,
	dataout_h_0,
	mac_rx_clock_connection_clk,
	mac_rgmii_connection_rx_control)/* synthesis synthesis_greybox=1 */;
output 	dataout_l_0;
output 	dataout_h_0;
input 	mac_rx_clock_connection_clk;
input 	mac_rgmii_connection_rx_control;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altddio_in_1 altddio_in_component(
	.dataout_l({dataout_l_unconnected_wire_3,dataout_l_unconnected_wire_2,dataout_l_unconnected_wire_1,dataout_l_0}),
	.dataout_h({dataout_h_unconnected_wire_3,dataout_h_unconnected_wire_2,dataout_h_unconnected_wire_1,dataout_h_0}),
	.inclock(mac_rx_clock_connection_clk),
	.datain({gnd,gnd,gnd,mac_rgmii_connection_rx_control}));

endmodule

module IoTOctopus_QSYS_altddio_in_1 (
	dataout_l,
	dataout_h,
	inclock,
	datain)/* synthesis synthesis_greybox=1 */;
output 	[3:0] dataout_l;
output 	[3:0] dataout_h;
input 	inclock;
input 	[3:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_ddio_in_gsd auto_generated(
	.dataout_l({dataout_l[0]}),
	.dataout_h({dataout_h[0]}),
	.inclock(inclock),
	.datain({datain[0]}));

endmodule

module IoTOctopus_QSYS_ddio_in_gsd (
	dataout_l,
	dataout_h,
	inclock,
	datain)/* synthesis synthesis_greybox=1 */;
output 	[0:0] dataout_l;
output 	[0:0] dataout_h;
input 	inclock;
input 	[0:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_in \ddio_ina[0] (
	.datain(datain[0]),
	.clk(inclock),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(dataout_l[0]),
	.regouthi(dataout_h[0]),
	.dfflo());
defparam \ddio_ina[0] .async_mode = "clear";
defparam \ddio_ina[0] .power_up = "low";
defparam \ddio_ina[0] .sync_mode = "none";
defparam \ddio_ina[0] .use_clkn = "false";

endmodule

module IoTOctopus_QSYS_altera_tse_rgmii_in4 (
	dataout_l_3,
	dataout_h_3,
	dataout_l_2,
	dataout_h_2,
	dataout_l_1,
	dataout_h_1,
	dataout_l_0,
	dataout_h_0,
	mac_rx_clock_connection_clk,
	mac_rgmii_connection_rgmii_in_3,
	mac_rgmii_connection_rgmii_in_2,
	mac_rgmii_connection_rgmii_in_1,
	mac_rgmii_connection_rgmii_in_0)/* synthesis synthesis_greybox=1 */;
output 	dataout_l_3;
output 	dataout_h_3;
output 	dataout_l_2;
output 	dataout_h_2;
output 	dataout_l_1;
output 	dataout_h_1;
output 	dataout_l_0;
output 	dataout_h_0;
input 	mac_rx_clock_connection_clk;
input 	mac_rgmii_connection_rgmii_in_3;
input 	mac_rgmii_connection_rgmii_in_2;
input 	mac_rgmii_connection_rgmii_in_1;
input 	mac_rgmii_connection_rgmii_in_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altddio_in_2 altddio_in_component(
	.dataout_l({dataout_l_3,dataout_l_2,dataout_l_1,dataout_l_0}),
	.dataout_h({dataout_h_3,dataout_h_2,dataout_h_1,dataout_h_0}),
	.inclock(mac_rx_clock_connection_clk),
	.datain({mac_rgmii_connection_rgmii_in_3,mac_rgmii_connection_rgmii_in_2,mac_rgmii_connection_rgmii_in_1,mac_rgmii_connection_rgmii_in_0}));

endmodule

module IoTOctopus_QSYS_altddio_in_2 (
	dataout_l,
	dataout_h,
	inclock,
	datain)/* synthesis synthesis_greybox=1 */;
output 	[3:0] dataout_l;
output 	[3:0] dataout_h;
input 	inclock;
input 	[3:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_ddio_in_jsd auto_generated(
	.dataout_l({dataout_l[3],dataout_l[2],dataout_l[1],dataout_l[0]}),
	.dataout_h({dataout_h[3],dataout_h[2],dataout_h[1],dataout_h[0]}),
	.inclock(inclock),
	.datain({datain[3],datain[2],datain[1],datain[0]}));

endmodule

module IoTOctopus_QSYS_ddio_in_jsd (
	dataout_l,
	dataout_h,
	inclock,
	datain)/* synthesis synthesis_greybox=1 */;
output 	[3:0] dataout_l;
output 	[3:0] dataout_h;
input 	inclock;
input 	[3:0] datain;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_in \ddio_ina[3] (
	.datain(datain[3]),
	.clk(inclock),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(dataout_l[3]),
	.regouthi(dataout_h[3]),
	.dfflo());
defparam \ddio_ina[3] .async_mode = "clear";
defparam \ddio_ina[3] .power_up = "low";
defparam \ddio_ina[3] .sync_mode = "none";
defparam \ddio_ina[3] .use_clkn = "false";

cyclonev_ddio_in \ddio_ina[2] (
	.datain(datain[2]),
	.clk(inclock),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(dataout_l[2]),
	.regouthi(dataout_h[2]),
	.dfflo());
defparam \ddio_ina[2] .async_mode = "clear";
defparam \ddio_ina[2] .power_up = "low";
defparam \ddio_ina[2] .sync_mode = "none";
defparam \ddio_ina[2] .use_clkn = "false";

cyclonev_ddio_in \ddio_ina[1] (
	.datain(datain[1]),
	.clk(inclock),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(dataout_l[1]),
	.regouthi(dataout_h[1]),
	.dfflo());
defparam \ddio_ina[1] .async_mode = "clear";
defparam \ddio_ina[1] .power_up = "low";
defparam \ddio_ina[1] .sync_mode = "none";
defparam \ddio_ina[1] .use_clkn = "false";

cyclonev_ddio_in \ddio_ina[0] (
	.datain(datain[0]),
	.clk(inclock),
	.clkn(gnd),
	.ena(vcc),
	.areset(gnd),
	.sreset(gnd),
	.regoutlo(dataout_l[0]),
	.regouthi(dataout_h[0]),
	.dfflo());
defparam \ddio_ina[0] .async_mode = "clear";
defparam \ddio_ina[0] .power_up = "low";
defparam \ddio_ina[0] .sync_mode = "none";
defparam \ddio_ina[0] .use_clkn = "false";

endmodule

module IoTOctopus_QSYS_altera_tse_rgmii_out1 (
	dataout_0,
	altera_tse_reset_synchronizer_chain_out,
	rgmii_out_1_wire_inp2,
	rgmii_out_1_wire_inp1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dataout_0;
input 	altera_tse_reset_synchronizer_chain_out;
input 	rgmii_out_1_wire_inp2;
input 	rgmii_out_1_wire_inp1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altddio_out_1 altddio_out_component(
	.dataout({gnd,gnd,gnd,dataout_0}),
	.aclr(altera_tse_reset_synchronizer_chain_out),
	.datain_l({gnd,gnd,gnd,rgmii_out_1_wire_inp2}),
	.datain_h({gnd,gnd,gnd,rgmii_out_1_wire_inp1}),
	.outclock(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altddio_out_1 (
	dataout,
	aclr,
	datain_l,
	datain_h,
	outclock)/* synthesis synthesis_greybox=1 */;
inout 	[3:0] dataout;
input 	aclr;
input 	[3:0] datain_l;
input 	[3:0] datain_h;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_ddio_out_ghb auto_generated(
	.dataout({dataout[0]}),
	.aclr(aclr),
	.datain_l({datain_l[0]}),
	.datain_h({datain_h[0]}),
	.outclock(outclock));

endmodule

module IoTOctopus_QSYS_ddio_out_ghb (
	dataout,
	aclr,
	datain_l,
	datain_h,
	outclock)/* synthesis synthesis_greybox=1 */;
output 	[0:0] dataout;
input 	aclr;
input 	[0:0] datain_l;
input 	[0:0] datain_h;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

endmodule

module IoTOctopus_QSYS_altera_tse_rgmii_out4 (
	dataout_0,
	dataout_1,
	dataout_2,
	dataout_3,
	altera_tse_reset_synchronizer_chain_out,
	rgmii_out_4_wire_4,
	rgmii_out_4_wire_0,
	rgmii_out_4_wire_5,
	rgmii_out_4_wire_1,
	rgmii_out_4_wire_6,
	rgmii_out_4_wire_2,
	rgmii_out_4_wire_7,
	rgmii_out_4_wire_3,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dataout_0;
output 	dataout_1;
output 	dataout_2;
output 	dataout_3;
input 	altera_tse_reset_synchronizer_chain_out;
input 	rgmii_out_4_wire_4;
input 	rgmii_out_4_wire_0;
input 	rgmii_out_4_wire_5;
input 	rgmii_out_4_wire_1;
input 	rgmii_out_4_wire_6;
input 	rgmii_out_4_wire_2;
input 	rgmii_out_4_wire_7;
input 	rgmii_out_4_wire_3;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altddio_out_2 altddio_out_component(
	.dataout({dataout_3,dataout_2,dataout_1,dataout_0}),
	.aclr(altera_tse_reset_synchronizer_chain_out),
	.datain_l({rgmii_out_4_wire_7,rgmii_out_4_wire_6,rgmii_out_4_wire_5,rgmii_out_4_wire_4}),
	.datain_h({rgmii_out_4_wire_3,rgmii_out_4_wire_2,rgmii_out_4_wire_1,rgmii_out_4_wire_0}),
	.outclock(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altddio_out_2 (
	dataout,
	aclr,
	datain_l,
	datain_h,
	outclock)/* synthesis synthesis_greybox=1 */;
inout 	[3:0] dataout;
input 	aclr;
input 	[3:0] datain_l;
input 	[3:0] datain_h;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_ddio_out_jhb auto_generated(
	.dataout({dataout[3],dataout[2],dataout[1],dataout[0]}),
	.aclr(aclr),
	.datain_l({datain_l[3],datain_l[2],datain_l[1],datain_l[0]}),
	.datain_h({datain_h[3],datain_h[2],datain_h[1],datain_h[0]}),
	.outclock(outclock));

endmodule

module IoTOctopus_QSYS_ddio_out_jhb (
	dataout,
	aclr,
	datain_l,
	datain_h,
	outclock)/* synthesis synthesis_greybox=1 */;
output 	[3:0] dataout;
input 	aclr;
input 	[3:0] datain_l;
input 	[3:0] datain_h;
input 	outclock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_ddio_out \ddio_outa[0] (
	.datainlo(datain_l[0]),
	.datainhi(datain_h[0]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[0]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[0] .async_mode = "clear";
defparam \ddio_outa[0] .half_rate_mode = "false";
defparam \ddio_outa[0] .power_up = "low";
defparam \ddio_outa[0] .sync_mode = "none";
defparam \ddio_outa[0] .use_new_clocking_model = "true";

cyclonev_ddio_out \ddio_outa[1] (
	.datainlo(datain_l[1]),
	.datainhi(datain_h[1]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[1]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[1] .async_mode = "clear";
defparam \ddio_outa[1] .half_rate_mode = "false";
defparam \ddio_outa[1] .power_up = "low";
defparam \ddio_outa[1] .sync_mode = "none";
defparam \ddio_outa[1] .use_new_clocking_model = "true";

cyclonev_ddio_out \ddio_outa[2] (
	.datainlo(datain_l[2]),
	.datainhi(datain_h[2]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[2]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[2] .async_mode = "clear";
defparam \ddio_outa[2] .half_rate_mode = "false";
defparam \ddio_outa[2] .power_up = "low";
defparam \ddio_outa[2] .sync_mode = "none";
defparam \ddio_outa[2] .use_new_clocking_model = "true";

cyclonev_ddio_out \ddio_outa[3] (
	.datainlo(datain_l[3]),
	.datainhi(datain_h[3]),
	.clkhi(outclock),
	.clklo(outclock),
	.muxsel(outclock),
	.ena(vcc),
	.areset(!aclr),
	.sreset(gnd),
	.hrbypass(gnd),
	.clk(gnd),
	.dataout(dataout[3]),
	.dfflo(),
	.dffhi());
defparam \ddio_outa[3] .async_mode = "clear";
defparam \ddio_outa[3] .half_rate_mode = "false";
defparam \ddio_outa[3] .power_up = "low";
defparam \ddio_outa[3] .sync_mode = "none";
defparam \ddio_outa[3] .use_new_clocking_model = "true";

endmodule

module IoTOctopus_QSYS_altera_tse_top_mdio (
	mdio_clk,
	mdio_out1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	mdio_clk;
output 	mdio_out1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mdio_out_int_reg1~q ;


IoTOctopus_QSYS_altera_tse_mdio_clk_gen U_CLKGEN(
	.mdio_clk1(mdio_clk),
	.reset(altera_tse_reset_synchronizer_chain_out),
	.reg_clk(clk_32_clk));

dffeas mdio_out(
	.clk(clk_32_clk),
	.d(\mdio_out_int_reg1~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mdio_out1),
	.prn(vcc));
defparam mdio_out.is_wysiwyg = "true";
defparam mdio_out.power_up = "low";

dffeas mdio_out_int_reg1(
	.clk(clk_32_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mdio_out_int_reg1~q ),
	.prn(vcc));
defparam mdio_out_int_reg1.is_wysiwyg = "true";
defparam mdio_out_int_reg1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_mdio_clk_gen (
	mdio_clk1,
	reset,
	reg_clk)/* synthesis synthesis_greybox=1 */;
output 	mdio_clk1;
input 	reset;
input 	reg_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~29_sumout ;
wire \Add0~2 ;
wire \Add0~21_sumout ;
wire \cnt[6]~q ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \cnt[7]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \cnt[0]~q ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \cnt[1]~q ;
wire \Add0~26 ;
wire \Add0~13_sumout ;
wire \cnt[2]~q ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \cnt[3]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \cnt[4]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \cnt[5]~q ;
wire \LessThan0~0_combout ;


dffeas mdio_clk(
	.clk(reg_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mdio_clk1),
	.prn(vcc));
defparam mdio_clk.is_wysiwyg = "true";
defparam mdio_clk.power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \cnt[6] (
	.clk(reg_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[6]~q ),
	.prn(vcc));
defparam \cnt[6] .is_wysiwyg = "true";
defparam \cnt[6] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \cnt[7] (
	.clk(reg_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[7]~q ),
	.prn(vcc));
defparam \cnt[7] .is_wysiwyg = "true";
defparam \cnt[7] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\cnt[5]~q ),
	.datab(!\cnt[4]~q ),
	.datac(!\cnt[1]~q ),
	.datad(!\cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\cnt[3]~q ),
	.datab(!\cnt[2]~q ),
	.datac(!\cnt[7]~q ),
	.datad(!\cnt[6]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \Equal0~1 .shared_arith = "off";

dffeas \cnt[0] (
	.clk(reg_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[0]~q ),
	.prn(vcc));
defparam \cnt[0] .is_wysiwyg = "true";
defparam \cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \cnt[1] (
	.clk(reg_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[1]~q ),
	.prn(vcc));
defparam \cnt[1] .is_wysiwyg = "true";
defparam \cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \cnt[2] (
	.clk(reg_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[2]~q ),
	.prn(vcc));
defparam \cnt[2] .is_wysiwyg = "true";
defparam \cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \cnt[3] (
	.clk(reg_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[3]~q ),
	.prn(vcc));
defparam \cnt[3] .is_wysiwyg = "true";
defparam \cnt[3] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \cnt[4] (
	.clk(reg_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[4]~q ),
	.prn(vcc));
defparam \cnt[4] .is_wysiwyg = "true";
defparam \cnt[4] .power_up = "low";

dffeas \cnt[5] (
	.clk(reg_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal0~1_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\cnt[5]~q ),
	.prn(vcc));
defparam \cnt[5] .is_wysiwyg = "true";
defparam \cnt[5] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\cnt[5]~q ),
	.datab(!\cnt[4]~q ),
	.datac(!\cnt[3]~q ),
	.datad(!\cnt[2]~q ),
	.datae(!\cnt[7]~q ),
	.dataf(!\cnt[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_top_w_fifo_10_100_1000 (
	gm_tx_d_reg_4,
	gm_tx_d_reg_0,
	gm_tx_d_reg_5,
	gm_tx_d_reg_1,
	gm_tx_d_reg_6,
	gm_tx_d_reg_2,
	gm_tx_d_reg_7,
	gm_tx_d_reg_3,
	gm_tx_err_reg,
	gm_tx_en_reg,
	septy_flag,
	tx_ff_uflow,
	afull_flag,
	aempty_flag,
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	ff_rx_err_stat_5,
	ff_rx_err_stat_6,
	ff_rx_err_stat_7,
	ff_rx_err_stat_8,
	ff_rx_err_stat_9,
	ff_rx_err_stat_10,
	ff_rx_err_stat_11,
	ff_rx_err_stat_12,
	ff_rx_err_stat_13,
	ff_rx_err_stat_14,
	ff_rx_err_stat_15,
	ff_rx_err_stat_16,
	ff_rx_err_stat_17,
	ff_rx_err_stat_18,
	ff_rx_err_stat_19,
	ff_rx_err_stat_20,
	ff_rx_err_stat_4,
	ff_rx_err_stat_22,
	ff_rx_ucast,
	ff_rx_mcast,
	ff_rx_bcast,
	ff_rx_vlan,
	sav_flag,
	afull_flag1,
	aempty_flag1,
	altera_tse_reset_synchronizer_chain_out,
	altera_tse_reset_synchronizer_chain_out1,
	altera_tse_reset_synchronizer_chain_out2,
	altera_tse_reset_synchronizer_chain_out3,
	mii_txd_int_0,
	mii_txd_int_1,
	mii_txd_int_2,
	mii_txd_int_3,
	mii_txerr_int,
	mii_txdv_int,
	LessThan0,
	magic_detect,
	ethernet_mode,
	sleep_ena,
	dreg_1,
	rx_dv,
	rgmii_in_4_reg_7,
	rgmii_in_4_reg_6,
	rgmii_in_4_reg_5,
	rgmii_in_4_reg_4,
	rgmii_in_4_reg_0,
	rgmii_in_4_reg_3,
	rgmii_in_4_reg_2,
	rgmii_in_4_reg_1,
	m_rx_crs,
	neinyesfmd,
	gm_rx_err,
	din_s1,
	GND_port,
	NJQG9082,
	clk_32_clk,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk,
	mac_misc_connection_ff_tx_crc_fwd)/* synthesis synthesis_greybox=1 */;
output 	gm_tx_d_reg_4;
output 	gm_tx_d_reg_0;
output 	gm_tx_d_reg_5;
output 	gm_tx_d_reg_1;
output 	gm_tx_d_reg_6;
output 	gm_tx_d_reg_2;
output 	gm_tx_d_reg_7;
output 	gm_tx_d_reg_3;
output 	gm_tx_err_reg;
output 	gm_tx_en_reg;
output 	septy_flag;
output 	tx_ff_uflow;
output 	afull_flag;
output 	aempty_flag;
output 	stateLOC_STATE_DATA;
output 	stateLOC_STATE_SHIFT;
output 	ff_rx_err_stat_5;
output 	ff_rx_err_stat_6;
output 	ff_rx_err_stat_7;
output 	ff_rx_err_stat_8;
output 	ff_rx_err_stat_9;
output 	ff_rx_err_stat_10;
output 	ff_rx_err_stat_11;
output 	ff_rx_err_stat_12;
output 	ff_rx_err_stat_13;
output 	ff_rx_err_stat_14;
output 	ff_rx_err_stat_15;
output 	ff_rx_err_stat_16;
output 	ff_rx_err_stat_17;
output 	ff_rx_err_stat_18;
output 	ff_rx_err_stat_19;
output 	ff_rx_err_stat_20;
output 	ff_rx_err_stat_4;
output 	ff_rx_err_stat_22;
output 	ff_rx_ucast;
output 	ff_rx_mcast;
output 	ff_rx_bcast;
output 	ff_rx_vlan;
output 	sav_flag;
output 	afull_flag1;
output 	aempty_flag1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_tse_reset_synchronizer_chain_out2;
input 	altera_tse_reset_synchronizer_chain_out3;
output 	mii_txd_int_0;
output 	mii_txd_int_1;
output 	mii_txd_int_2;
output 	mii_txd_int_3;
output 	mii_txerr_int;
output 	mii_txdv_int;
input 	LessThan0;
output 	magic_detect;
input 	ethernet_mode;
input 	sleep_ena;
input 	dreg_1;
input 	rx_dv;
input 	rgmii_in_4_reg_7;
input 	rgmii_in_4_reg_6;
input 	rgmii_in_4_reg_5;
input 	rgmii_in_4_reg_4;
input 	rgmii_in_4_reg_0;
input 	rgmii_in_4_reg_3;
input 	rgmii_in_4_reg_2;
input 	rgmii_in_4_reg_1;
input 	m_rx_crs;
output 	neinyesfmd;
input 	gm_rx_err;
output 	din_s1;
input 	GND_port;
input 	NJQG9082;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;
input 	mac_misc_connection_ff_tx_crc_fwd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_LBFF|en~q ;
wire \U_LBFF|data[3]~q ;
wire \U_LBFF|data[2]~q ;
wire \U_LBFF|data[1]~q ;
wire \U_LBFF|data[0]~q ;
wire \U_LBFF|data[7]~q ;
wire \U_LBFF|data[6]~q ;
wire \U_LBFF|data[5]~q ;
wire \U_LBFF|data[4]~q ;
wire \U_MRX|mii_rxd_o[3]~q ;
wire \U_MRX|mii_rxd_o[2]~q ;
wire \U_MRX|mii_rxd_o[1]~q ;
wire \U_MRX|mii_rxd_o[0]~q ;
wire \U_MRX|mii_rxd_o[7]~q ;
wire \U_MRX|mii_rxd_o[6]~q ;
wire \U_MRX|mii_rxd_o[5]~q ;
wire \U_MRX|mii_rxd_o[4]~q ;
wire \U_LBFF|err~q ;
wire \U_MRX|mii_rxerr_o~q ;
wire \U_CLKCT|txclk_ena~q ;
wire \U_MAC|U_GETH|U_TX|tx_en_s[1]~q ;
wire \U_CLKCT|rxclk_ena~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[4]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[0]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[5]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[1]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[6]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[2]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[7]~q ;
wire \U_MAC|U_GETH|U_TX|rd_14[3]~q ;
wire \U_MAC|U_GETH|U_TX|tx_err~q ;
wire \U_MRX|mii_clk_ena~q ;
wire \U_SYNC_2|std_sync_no_cut|dreg[1]~q ;
wire \U_GMIF|gm_rx_en_i_reg~q ;
wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \U_MRX|packet_in_progress~q ;
wire \U_GMIF|gm_rx_d_i_reg[3]~q ;
wire \U_GMIF|gm_rx_d_i_reg[2]~q ;
wire \U_GMIF|gm_rx_d_i_reg[1]~q ;
wire \U_GMIF|gm_rx_d_i_reg[0]~q ;
wire \U_GMIF|gm_rx_d_i_reg[7]~q ;
wire \U_GMIF|gm_rx_d_i_reg[6]~q ;
wire \U_GMIF|gm_rx_d_i_reg[5]~q ;
wire \U_GMIF|gm_rx_d_i_reg[4]~q ;
wire \U_GMIF|gm_rx_err_i_reg~q ;


IoTOctopus_QSYS_altera_tse_top_w_fifo U_MAC(
	.en(\U_LBFF|en~q ),
	.data_3(\U_LBFF|data[3]~q ),
	.data_2(\U_LBFF|data[2]~q ),
	.data_1(\U_LBFF|data[1]~q ),
	.data_0(\U_LBFF|data[0]~q ),
	.data_7(\U_LBFF|data[7]~q ),
	.data_6(\U_LBFF|data[6]~q ),
	.data_5(\U_LBFF|data[5]~q ),
	.data_4(\U_LBFF|data[4]~q ),
	.err(\U_LBFF|err~q ),
	.septy_flag(septy_flag),
	.tx_ff_uflow(tx_ff_uflow),
	.afull_flag(afull_flag),
	.aempty_flag(aempty_flag),
	.stateLOC_STATE_DATA(stateLOC_STATE_DATA),
	.stateLOC_STATE_SHIFT(stateLOC_STATE_SHIFT),
	.ff_rx_err_stat_5(ff_rx_err_stat_5),
	.ff_rx_err_stat_6(ff_rx_err_stat_6),
	.ff_rx_err_stat_7(ff_rx_err_stat_7),
	.ff_rx_err_stat_8(ff_rx_err_stat_8),
	.ff_rx_err_stat_9(ff_rx_err_stat_9),
	.ff_rx_err_stat_10(ff_rx_err_stat_10),
	.ff_rx_err_stat_11(ff_rx_err_stat_11),
	.ff_rx_err_stat_12(ff_rx_err_stat_12),
	.ff_rx_err_stat_13(ff_rx_err_stat_13),
	.ff_rx_err_stat_14(ff_rx_err_stat_14),
	.ff_rx_err_stat_15(ff_rx_err_stat_15),
	.ff_rx_err_stat_16(ff_rx_err_stat_16),
	.ff_rx_err_stat_17(ff_rx_err_stat_17),
	.ff_rx_err_stat_18(ff_rx_err_stat_18),
	.ff_rx_err_stat_19(ff_rx_err_stat_19),
	.ff_rx_err_stat_20(ff_rx_err_stat_20),
	.ff_rx_err_stat_4(ff_rx_err_stat_4),
	.ff_rx_err_stat_22(ff_rx_err_stat_22),
	.ff_rx_ucast(ff_rx_ucast),
	.ff_rx_mcast(ff_rx_mcast),
	.ff_rx_bcast(ff_rx_bcast),
	.ff_rx_vlan(ff_rx_vlan),
	.sav_flag(sav_flag),
	.afull_flag1(afull_flag1),
	.aempty_flag1(aempty_flag1),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.txclk_ena(\U_CLKCT|txclk_ena~q ),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.altera_tse_reset_synchronizer_chain_out2(altera_tse_reset_synchronizer_chain_out2),
	.altera_tse_reset_synchronizer_chain_out3(altera_tse_reset_synchronizer_chain_out3),
	.tx_en_s_1(\U_MAC|U_GETH|U_TX|tx_en_s[1]~q ),
	.rxclk_ena(\U_CLKCT|rxclk_ena~q ),
	.LessThan0(LessThan0),
	.rd_14_4(\U_MAC|U_GETH|U_TX|rd_14[4]~q ),
	.rd_14_0(\U_MAC|U_GETH|U_TX|rd_14[0]~q ),
	.rd_14_5(\U_MAC|U_GETH|U_TX|rd_14[5]~q ),
	.rd_14_1(\U_MAC|U_GETH|U_TX|rd_14[1]~q ),
	.rd_14_6(\U_MAC|U_GETH|U_TX|rd_14[6]~q ),
	.rd_14_2(\U_MAC|U_GETH|U_TX|rd_14[2]~q ),
	.rd_14_7(\U_MAC|U_GETH|U_TX|rd_14[7]~q ),
	.rd_14_3(\U_MAC|U_GETH|U_TX|rd_14[3]~q ),
	.tx_err(\U_MAC|U_GETH|U_TX|tx_err~q ),
	.magic_detect(magic_detect),
	.ethernet_mode(ethernet_mode),
	.sleep_ena(sleep_ena),
	.dreg_1(dreg_1),
	.m_rx_crs(m_rx_crs),
	.dreg_11(\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.din_s1(din_s1),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk),
	.mac_misc_connection_ff_tx_crc_fwd(mac_misc_connection_ff_tx_crc_fwd));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_17 U_SYNC_2(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_loopback_ff U_LBFF(
	.en1(\U_LBFF|en~q ),
	.data_3(\U_LBFF|data[3]~q ),
	.data_2(\U_LBFF|data[2]~q ),
	.data_1(\U_LBFF|data[1]~q ),
	.data_0(\U_LBFF|data[0]~q ),
	.data_7(\U_LBFF|data[7]~q ),
	.data_6(\U_LBFF|data[6]~q ),
	.data_5(\U_LBFF|data[5]~q ),
	.data_4(\U_LBFF|data[4]~q ),
	.mii_rxd_o_3(\U_MRX|mii_rxd_o[3]~q ),
	.mii_rxd_o_2(\U_MRX|mii_rxd_o[2]~q ),
	.mii_rxd_o_1(\U_MRX|mii_rxd_o[1]~q ),
	.mii_rxd_o_0(\U_MRX|mii_rxd_o[0]~q ),
	.mii_rxd_o_7(\U_MRX|mii_rxd_o[7]~q ),
	.mii_rxd_o_6(\U_MRX|mii_rxd_o[6]~q ),
	.mii_rxd_o_5(\U_MRX|mii_rxd_o[5]~q ),
	.mii_rxd_o_4(\U_MRX|mii_rxd_o[4]~q ),
	.err1(\U_LBFF|err~q ),
	.mii_rxerr_o(\U_MRX|mii_rxerr_o~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out3),
	.tx_en_s_1(\U_MAC|U_GETH|U_TX|tx_en_s[1]~q ),
	.rd_14_4(\U_MAC|U_GETH|U_TX|rd_14[4]~q ),
	.rd_14_0(\U_MAC|U_GETH|U_TX|rd_14[0]~q ),
	.rd_14_5(\U_MAC|U_GETH|U_TX|rd_14[5]~q ),
	.rd_14_1(\U_MAC|U_GETH|U_TX|rd_14[1]~q ),
	.rd_14_6(\U_MAC|U_GETH|U_TX|rd_14[6]~q ),
	.rd_14_2(\U_MAC|U_GETH|U_TX|rd_14[2]~q ),
	.rd_14_7(\U_MAC|U_GETH|U_TX|rd_14[7]~q ),
	.rd_14_3(\U_MAC|U_GETH|U_TX|rd_14[3]~q ),
	.tx_err(\U_MAC|U_GETH|U_TX|tx_err~q ),
	.gm_rx_en_i_reg(\U_GMIF|gm_rx_en_i_reg~q ),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.packet_in_progress(\U_MRX|packet_in_progress~q ),
	.gm_rx_d_i_reg_3(\U_GMIF|gm_rx_d_i_reg[3]~q ),
	.gm_rx_d_i_reg_2(\U_GMIF|gm_rx_d_i_reg[2]~q ),
	.gm_rx_d_i_reg_1(\U_GMIF|gm_rx_d_i_reg[1]~q ),
	.gm_rx_d_i_reg_0(\U_GMIF|gm_rx_d_i_reg[0]~q ),
	.gm_rx_d_i_reg_7(\U_GMIF|gm_rx_d_i_reg[7]~q ),
	.gm_rx_d_i_reg_6(\U_GMIF|gm_rx_d_i_reg[6]~q ),
	.gm_rx_d_i_reg_5(\U_GMIF|gm_rx_d_i_reg[5]~q ),
	.gm_rx_d_i_reg_4(\U_GMIF|gm_rx_d_i_reg[4]~q ),
	.gm_rx_err_i_reg(\U_GMIF|gm_rx_err_i_reg~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_16 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out3),
	.ethernet_mode(ethernet_mode),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gmii_io U_GMIF(
	.gm_tx_d_reg_4(gm_tx_d_reg_4),
	.gm_tx_d_reg_0(gm_tx_d_reg_0),
	.gm_tx_d_reg_5(gm_tx_d_reg_5),
	.gm_tx_d_reg_1(gm_tx_d_reg_1),
	.gm_tx_d_reg_6(gm_tx_d_reg_6),
	.gm_tx_d_reg_2(gm_tx_d_reg_2),
	.gm_tx_d_reg_7(gm_tx_d_reg_7),
	.gm_tx_d_reg_3(gm_tx_d_reg_3),
	.gm_tx_err_reg1(gm_tx_err_reg),
	.gm_tx_en_reg1(gm_tx_en_reg),
	.reset_tx_clk(altera_tse_reset_synchronizer_chain_out1),
	.reset_rx_clk(altera_tse_reset_synchronizer_chain_out3),
	.tx_en_s_1(\U_MAC|U_GETH|U_TX|tx_en_s[1]~q ),
	.rd_14_4(\U_MAC|U_GETH|U_TX|rd_14[4]~q ),
	.rd_14_0(\U_MAC|U_GETH|U_TX|rd_14[0]~q ),
	.rd_14_5(\U_MAC|U_GETH|U_TX|rd_14[5]~q ),
	.rd_14_1(\U_MAC|U_GETH|U_TX|rd_14[1]~q ),
	.rd_14_6(\U_MAC|U_GETH|U_TX|rd_14[6]~q ),
	.rd_14_2(\U_MAC|U_GETH|U_TX|rd_14[2]~q ),
	.rd_14_7(\U_MAC|U_GETH|U_TX|rd_14[7]~q ),
	.rd_14_3(\U_MAC|U_GETH|U_TX|rd_14[3]~q ),
	.tx_err(\U_MAC|U_GETH|U_TX|tx_err~q ),
	.ethernet_mode(ethernet_mode),
	.gm_rx_en(rx_dv),
	.gm_rx_d({rgmii_in_4_reg_7,rgmii_in_4_reg_6,rgmii_in_4_reg_5,rgmii_in_4_reg_4,rgmii_in_4_reg_3,rgmii_in_4_reg_2,rgmii_in_4_reg_1,rgmii_in_4_reg_0}),
	.gm_rx_en_i_reg1(\U_GMIF|gm_rx_en_i_reg~q ),
	.gm_rx_d_i_reg_3(\U_GMIF|gm_rx_d_i_reg[3]~q ),
	.gm_rx_d_i_reg_2(\U_GMIF|gm_rx_d_i_reg[2]~q ),
	.gm_rx_d_i_reg_1(\U_GMIF|gm_rx_d_i_reg[1]~q ),
	.gm_rx_d_i_reg_0(\U_GMIF|gm_rx_d_i_reg[0]~q ),
	.gm_rx_d_i_reg_7(\U_GMIF|gm_rx_d_i_reg[7]~q ),
	.gm_rx_d_i_reg_6(\U_GMIF|gm_rx_d_i_reg[6]~q ),
	.gm_rx_d_i_reg_5(\U_GMIF|gm_rx_d_i_reg[5]~q ),
	.gm_rx_d_i_reg_4(\U_GMIF|gm_rx_d_i_reg[4]~q ),
	.gm_rx_err_i_reg1(\U_GMIF|gm_rx_err_i_reg~q ),
	.gm_rx_err(gm_rx_err),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.rx_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_mii_tx_if U_MTX(
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.mii_txd_int_0(mii_txd_int_0),
	.mii_txd_int_1(mii_txd_int_1),
	.mii_txd_int_2(mii_txd_int_2),
	.mii_txd_int_3(mii_txd_int_3),
	.mii_txerr_int1(mii_txerr_int),
	.mii_txdv_int1(mii_txdv_int),
	.tx_en_s_1(\U_MAC|U_GETH|U_TX|tx_en_s[1]~q ),
	.rd_14_4(\U_MAC|U_GETH|U_TX|rd_14[4]~q ),
	.rd_14_0(\U_MAC|U_GETH|U_TX|rd_14[0]~q ),
	.rd_14_5(\U_MAC|U_GETH|U_TX|rd_14[5]~q ),
	.rd_14_1(\U_MAC|U_GETH|U_TX|rd_14[1]~q ),
	.rd_14_6(\U_MAC|U_GETH|U_TX|rd_14[6]~q ),
	.rd_14_2(\U_MAC|U_GETH|U_TX|rd_14[2]~q ),
	.rd_14_7(\U_MAC|U_GETH|U_TX|rd_14[7]~q ),
	.rd_14_3(\U_MAC|U_GETH|U_TX|rd_14[3]~q ),
	.tx_err(\U_MAC|U_GETH|U_TX|tx_err~q ),
	.ethernet_mode(ethernet_mode),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_mii_rx_if U_MRX(
	.mii_rxd_o_3(\U_MRX|mii_rxd_o[3]~q ),
	.mii_rxd_o_2(\U_MRX|mii_rxd_o[2]~q ),
	.mii_rxd_o_1(\U_MRX|mii_rxd_o[1]~q ),
	.mii_rxd_o_0(\U_MRX|mii_rxd_o[0]~q ),
	.mii_rxd_o_7(\U_MRX|mii_rxd_o[7]~q ),
	.mii_rxd_o_6(\U_MRX|mii_rxd_o[6]~q ),
	.mii_rxd_o_5(\U_MRX|mii_rxd_o[5]~q ),
	.mii_rxd_o_4(\U_MRX|mii_rxd_o[4]~q ),
	.mii_rxerr_o1(\U_MRX|mii_rxerr_o~q ),
	.reset(altera_tse_reset_synchronizer_chain_out3),
	.mii_clk_ena1(\U_MRX|mii_clk_ena~q ),
	.gm_rx_en_i_reg(\U_GMIF|gm_rx_en_i_reg~q ),
	.packet_in_progress1(\U_MRX|packet_in_progress~q ),
	.gm_rx_d_i_reg_3(\U_GMIF|gm_rx_d_i_reg[3]~q ),
	.gm_rx_d_i_reg_2(\U_GMIF|gm_rx_d_i_reg[2]~q ),
	.gm_rx_d_i_reg_1(\U_GMIF|gm_rx_d_i_reg[1]~q ),
	.gm_rx_d_i_reg_0(\U_GMIF|gm_rx_d_i_reg[0]~q ),
	.gm_rx_err_i_reg(\U_GMIF|gm_rx_err_i_reg~q ),
	.rx_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_clk_cntl U_CLKCT(
	.txclk_ena1(\U_CLKCT|txclk_ena~q ),
	.reset_tx_clk(altera_tse_reset_synchronizer_chain_out1),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out3),
	.rxclk_ena1(\U_CLKCT|rxclk_ena~q ),
	.mii_clk_ena(\U_MRX|mii_clk_ena~q ),
	.ethernet_mode(ethernet_mode),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

cyclonev_lcell_comb \neinyesfmd~55 (
	.dataa(!NJQG9082),
	.datab(!mii_txdv_int),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(neinyesfmd),
	.sumout(),
	.cout(),
	.shareout());
defparam \neinyesfmd~55 .extended_lut = "off";
defparam \neinyesfmd~55 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \neinyesfmd~55 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_16 (
	altera_tse_reset_synchronizer_chain_out,
	ethernet_mode,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
input 	ethernet_mode;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_16 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.din(ethernet_mode),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_16 (
	reset_n,
	din,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_17 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_17 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_17 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_clk_cntl (
	txclk_ena1,
	reset_tx_clk,
	altera_tse_reset_synchronizer_chain_out,
	rxclk_ena1,
	mii_clk_ena,
	ethernet_mode,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	txclk_ena1;
input 	reset_tx_clk;
input 	altera_tse_reset_synchronizer_chain_out;
output 	rxclk_ena1;
input 	mii_clk_ena;
input 	ethernet_mode;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_TX_ETH_MODE|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_RX_ETH_MODE|std_sync_no_cut|dreg[1]~q ;
wire \txclk_ena_i~0_combout ;
wire \txclk_ena_i~q ;
wire \txclk_ena~0_combout ;
wire \rxclk_ena~0_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_19 U_SYNC_TX_ETH_MODE(
	.altera_tse_reset_synchronizer_chain_out(reset_tx_clk),
	.dreg_1(\U_SYNC_TX_ETH_MODE|std_sync_no_cut|dreg[1]~q ),
	.ethernet_mode(ethernet_mode),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_18 U_SYNC_RX_ETH_MODE(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_RX_ETH_MODE|std_sync_no_cut|dreg[1]~q ),
	.ethernet_mode(ethernet_mode),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

dffeas txclk_ena(
	.clk(mac_tx_clock_connection_clk),
	.d(\txclk_ena~0_combout ),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(txclk_ena1),
	.prn(vcc));
defparam txclk_ena.is_wysiwyg = "true";
defparam txclk_ena.power_up = "low";

dffeas rxclk_ena(
	.clk(mac_rx_clock_connection_clk),
	.d(\rxclk_ena~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rxclk_ena1),
	.prn(vcc));
defparam rxclk_ena.is_wysiwyg = "true";
defparam rxclk_ena.power_up = "low";

cyclonev_lcell_comb \txclk_ena_i~0 (
	.dataa(!\txclk_ena_i~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\txclk_ena_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \txclk_ena_i~0 .extended_lut = "off";
defparam \txclk_ena_i~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \txclk_ena_i~0 .shared_arith = "off";

dffeas txclk_ena_i(
	.clk(mac_tx_clock_connection_clk),
	.d(\txclk_ena_i~0_combout ),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\txclk_ena_i~q ),
	.prn(vcc));
defparam txclk_ena_i.is_wysiwyg = "true";
defparam txclk_ena_i.power_up = "low";

cyclonev_lcell_comb \txclk_ena~0 (
	.dataa(!\txclk_ena_i~q ),
	.datab(!\U_SYNC_TX_ETH_MODE|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\txclk_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \txclk_ena~0 .extended_lut = "off";
defparam \txclk_ena~0 .lut_mask = 64'h7777777777777777;
defparam \txclk_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \rxclk_ena~0 (
	.dataa(!\U_SYNC_RX_ETH_MODE|std_sync_no_cut|dreg[1]~q ),
	.datab(!mii_clk_ena),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxclk_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxclk_ena~0 .extended_lut = "off";
defparam \rxclk_ena~0 .lut_mask = 64'h7777777777777777;
defparam \rxclk_ena~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_18 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	ethernet_mode,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	ethernet_mode;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_18 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(ethernet_mode),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_18 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_19 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	ethernet_mode,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	ethernet_mode;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_19 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(ethernet_mode),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_19 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_gmii_io (
	gm_tx_d_reg_4,
	gm_tx_d_reg_0,
	gm_tx_d_reg_5,
	gm_tx_d_reg_1,
	gm_tx_d_reg_6,
	gm_tx_d_reg_2,
	gm_tx_d_reg_7,
	gm_tx_d_reg_3,
	gm_tx_err_reg1,
	gm_tx_en_reg1,
	reset_tx_clk,
	reset_rx_clk,
	tx_en_s_1,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	ethernet_mode,
	gm_rx_en,
	gm_rx_d,
	gm_rx_en_i_reg1,
	gm_rx_d_i_reg_3,
	gm_rx_d_i_reg_2,
	gm_rx_d_i_reg_1,
	gm_rx_d_i_reg_0,
	gm_rx_d_i_reg_7,
	gm_rx_d_i_reg_6,
	gm_rx_d_i_reg_5,
	gm_rx_d_i_reg_4,
	gm_rx_err_i_reg1,
	gm_rx_err,
	mac_tx_clock_connection_clk,
	rx_clk)/* synthesis synthesis_greybox=1 */;
output 	gm_tx_d_reg_4;
output 	gm_tx_d_reg_0;
output 	gm_tx_d_reg_5;
output 	gm_tx_d_reg_1;
output 	gm_tx_d_reg_6;
output 	gm_tx_d_reg_2;
output 	gm_tx_d_reg_7;
output 	gm_tx_d_reg_3;
output 	gm_tx_err_reg1;
output 	gm_tx_en_reg1;
input 	reset_tx_clk;
input 	reset_rx_clk;
input 	tx_en_s_1;
input 	rd_14_4;
input 	rd_14_0;
input 	rd_14_5;
input 	rd_14_1;
input 	rd_14_6;
input 	rd_14_2;
input 	rd_14_7;
input 	rd_14_3;
input 	tx_err;
input 	ethernet_mode;
input 	gm_rx_en;
input 	[7:0] gm_rx_d;
output 	gm_rx_en_i_reg1;
output 	gm_rx_d_i_reg_3;
output 	gm_rx_d_i_reg_2;
output 	gm_rx_d_i_reg_1;
output 	gm_rx_d_i_reg_0;
output 	gm_rx_d_i_reg_7;
output 	gm_rx_d_i_reg_6;
output 	gm_rx_d_i_reg_5;
output 	gm_rx_d_i_reg_4;
output 	gm_rx_err_i_reg1;
input 	gm_rx_err;
input 	mac_tx_clock_connection_clk;
input 	rx_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_20 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(reset_tx_clk),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.ethernet_mode(ethernet_mode),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

dffeas \gm_tx_d_reg[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_4),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_4),
	.prn(vcc));
defparam \gm_tx_d_reg[4] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[4] .power_up = "low";

dffeas \gm_tx_d_reg[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_0),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_0),
	.prn(vcc));
defparam \gm_tx_d_reg[0] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[0] .power_up = "low";

dffeas \gm_tx_d_reg[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_5),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_5),
	.prn(vcc));
defparam \gm_tx_d_reg[5] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[5] .power_up = "low";

dffeas \gm_tx_d_reg[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_1),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_1),
	.prn(vcc));
defparam \gm_tx_d_reg[1] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[1] .power_up = "low";

dffeas \gm_tx_d_reg[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_6),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_6),
	.prn(vcc));
defparam \gm_tx_d_reg[6] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[6] .power_up = "low";

dffeas \gm_tx_d_reg[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_2),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_2),
	.prn(vcc));
defparam \gm_tx_d_reg[2] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[2] .power_up = "low";

dffeas \gm_tx_d_reg[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_7),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_7),
	.prn(vcc));
defparam \gm_tx_d_reg[7] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[7] .power_up = "low";

dffeas \gm_tx_d_reg[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(rd_14_3),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_d_reg_3),
	.prn(vcc));
defparam \gm_tx_d_reg[3] .is_wysiwyg = "true";
defparam \gm_tx_d_reg[3] .power_up = "low";

dffeas gm_tx_err_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(tx_err),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_err_reg1),
	.prn(vcc));
defparam gm_tx_err_reg.is_wysiwyg = "true";
defparam gm_tx_err_reg.power_up = "low";

dffeas gm_tx_en_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(tx_en_s_1),
	.asdata(vcc),
	.clrn(reset_tx_clk),
	.aload(gnd),
	.sclr(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(gm_tx_en_reg1),
	.prn(vcc));
defparam gm_tx_en_reg.is_wysiwyg = "true";
defparam gm_tx_en_reg.power_up = "low";

dffeas gm_rx_en_i_reg(
	.clk(rx_clk),
	.d(gm_rx_en),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_en_i_reg1),
	.prn(vcc));
defparam gm_rx_en_i_reg.is_wysiwyg = "true";
defparam gm_rx_en_i_reg.power_up = "low";

dffeas \gm_rx_d_i_reg[3] (
	.clk(rx_clk),
	.d(gm_rx_d[3]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_3),
	.prn(vcc));
defparam \gm_rx_d_i_reg[3] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[3] .power_up = "low";

dffeas \gm_rx_d_i_reg[2] (
	.clk(rx_clk),
	.d(gm_rx_d[2]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_2),
	.prn(vcc));
defparam \gm_rx_d_i_reg[2] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[2] .power_up = "low";

dffeas \gm_rx_d_i_reg[1] (
	.clk(rx_clk),
	.d(gm_rx_d[1]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_1),
	.prn(vcc));
defparam \gm_rx_d_i_reg[1] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[1] .power_up = "low";

dffeas \gm_rx_d_i_reg[0] (
	.clk(rx_clk),
	.d(gm_rx_d[0]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_0),
	.prn(vcc));
defparam \gm_rx_d_i_reg[0] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[0] .power_up = "low";

dffeas \gm_rx_d_i_reg[7] (
	.clk(rx_clk),
	.d(gm_rx_d[7]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_7),
	.prn(vcc));
defparam \gm_rx_d_i_reg[7] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[7] .power_up = "low";

dffeas \gm_rx_d_i_reg[6] (
	.clk(rx_clk),
	.d(gm_rx_d[6]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_6),
	.prn(vcc));
defparam \gm_rx_d_i_reg[6] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[6] .power_up = "low";

dffeas \gm_rx_d_i_reg[5] (
	.clk(rx_clk),
	.d(gm_rx_d[5]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_5),
	.prn(vcc));
defparam \gm_rx_d_i_reg[5] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[5] .power_up = "low";

dffeas \gm_rx_d_i_reg[4] (
	.clk(rx_clk),
	.d(gm_rx_d[4]),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_d_i_reg_4),
	.prn(vcc));
defparam \gm_rx_d_i_reg[4] .is_wysiwyg = "true";
defparam \gm_rx_d_i_reg[4] .power_up = "low";

dffeas gm_rx_err_i_reg(
	.clk(rx_clk),
	.d(gm_rx_err),
	.asdata(vcc),
	.clrn(reset_rx_clk),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(gm_rx_err_i_reg1),
	.prn(vcc));
defparam gm_rx_err_i_reg.is_wysiwyg = "true";
defparam gm_rx_err_i_reg.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_20 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	ethernet_mode,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	ethernet_mode;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_20 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(ethernet_mode),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_20 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_loopback_ff (
	en1,
	data_3,
	data_2,
	data_1,
	data_0,
	data_7,
	data_6,
	data_5,
	data_4,
	mii_rxd_o_3,
	mii_rxd_o_2,
	mii_rxd_o_1,
	mii_rxd_o_0,
	mii_rxd_o_7,
	mii_rxd_o_6,
	mii_rxd_o_5,
	mii_rxd_o_4,
	err1,
	mii_rxerr_o,
	altera_tse_reset_synchronizer_chain_out,
	altera_tse_reset_synchronizer_chain_out1,
	tx_en_s_1,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	gm_rx_en_i_reg,
	dreg_1,
	packet_in_progress,
	gm_rx_d_i_reg_3,
	gm_rx_d_i_reg_2,
	gm_rx_d_i_reg_1,
	gm_rx_d_i_reg_0,
	gm_rx_d_i_reg_7,
	gm_rx_d_i_reg_6,
	gm_rx_d_i_reg_5,
	gm_rx_d_i_reg_4,
	gm_rx_err_i_reg,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	en1;
output 	data_3;
output 	data_2;
output 	data_1;
output 	data_0;
output 	data_7;
output 	data_6;
output 	data_5;
output 	data_4;
input 	mii_rxd_o_3;
input 	mii_rxd_o_2;
input 	mii_rxd_o_1;
input 	mii_rxd_o_0;
input 	mii_rxd_o_7;
input 	mii_rxd_o_6;
input 	mii_rxd_o_5;
input 	mii_rxd_o_4;
output 	err1;
input 	mii_rxerr_o;
input 	altera_tse_reset_synchronizer_chain_out;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	tx_en_s_1;
input 	rd_14_4;
input 	rd_14_0;
input 	rd_14_5;
input 	rd_14_1;
input 	rd_14_6;
input 	rd_14_2;
input 	rd_14_7;
input 	rd_14_3;
input 	tx_err;
input 	gm_rx_en_i_reg;
input 	dreg_1;
input 	packet_in_progress;
input 	gm_rx_d_i_reg_3;
input 	gm_rx_d_i_reg_2;
input 	gm_rx_d_i_reg_1;
input 	gm_rx_d_i_reg_0;
input 	gm_rx_d_i_reg_7;
input 	gm_rx_d_i_reg_6;
input 	gm_rx_d_i_reg_5;
input 	gm_rx_d_i_reg_4;
input 	gm_rx_err_i_reg;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_LBR|ff_gmii_reg~q ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[8] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[3] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[2] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[1] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[0] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[7] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[6] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[5] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[4] ;
wire \U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[9] ;
wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \U_LBR|state.STM_TYPE_FRM_READ~q ;
wire \U_LBFF|aempty_flag~q ;
wire \U_LBR|state.STM_TYPE_IDLE~q ;
wire \U_LBR|Selector1~0_combout ;
wire \U_LBFF|aempty_low_det~q ;
wire \U_LBR|Selector1~1_combout ;
wire \U_LBFF|afull_flag~q ;
wire \U_LBW|ff_wren~0_combout ;
wire \en~0_combout ;
wire \data[7]~0_combout ;
wire \data_reg[3]~q ;
wire \data~1_combout ;
wire \data_reg[2]~q ;
wire \data~2_combout ;
wire \data_reg[1]~q ;
wire \data~3_combout ;
wire \data_reg[0]~q ;
wire \data~4_combout ;
wire \data_reg[7]~q ;
wire \data~5_combout ;
wire \data_reg[6]~q ;
wire \data~6_combout ;
wire \data_reg[5]~q ;
wire \data~7_combout ;
wire \data_reg[4]~q ;
wire \data~8_combout ;
wire \err_reg~q ;
wire \err~0_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_21 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_lb_read_cntl U_LBR(
	.ff_gmii_reg1(\U_LBR|ff_gmii_reg~q ),
	.ff_gmii_en(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[8] ),
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.stateSTM_TYPE_FRM_READ(\U_LBR|state.STM_TYPE_FRM_READ~q ),
	.aempty_flag(\U_LBFF|aempty_flag~q ),
	.stateSTM_TYPE_IDLE(\U_LBR|state.STM_TYPE_IDLE~q ),
	.Selector1(\U_LBR|Selector1~0_combout ),
	.aempty_low_det(\U_LBFF|aempty_low_det~q ),
	.Selector11(\U_LBR|Selector1~1_combout ),
	.clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_a_fifo_24 U_LBFF(
	.ff_gmii_reg(\U_LBR|ff_gmii_reg~q ),
	.q_b_8(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[8] ),
	.q_b_3(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.q_b_2(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.q_b_1(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.q_b_7(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[7] ),
	.q_b_6(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[6] ),
	.q_b_5(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[5] ),
	.q_b_4(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[4] ),
	.q_b_9(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[9] ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.tx_en_s_1(tx_en_s_1),
	.rd_14_4(rd_14_4),
	.rd_14_0(rd_14_0),
	.rd_14_5(rd_14_5),
	.rd_14_1(rd_14_1),
	.rd_14_6(rd_14_6),
	.rd_14_2(rd_14_2),
	.rd_14_7(rd_14_7),
	.rd_14_3(rd_14_3),
	.tx_err(tx_err),
	.stateSTM_TYPE_FRM_READ(\U_LBR|state.STM_TYPE_FRM_READ~q ),
	.aempty_flag1(\U_LBFF|aempty_flag~q ),
	.Selector1(\U_LBR|Selector1~0_combout ),
	.aempty_low_det1(\U_LBFF|aempty_low_det~q ),
	.Selector11(\U_LBR|Selector1~1_combout ),
	.afull_flag1(\U_LBFF|afull_flag~q ),
	.ff_wren(\U_LBW|ff_wren~0_combout ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_lb_wrt_cntl U_LBW(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.tx_en_s_1(tx_en_s_1),
	.afull_flag(\U_LBFF|afull_flag~q ),
	.ff_wren(\U_LBW|ff_wren~0_combout ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

dffeas en(
	.clk(mac_rx_clock_connection_clk),
	.d(\en~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(en1),
	.prn(vcc));
defparam en.is_wysiwyg = "true";
defparam en.power_up = "low";

dffeas \data[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_3),
	.prn(vcc));
defparam \data[3] .is_wysiwyg = "true";
defparam \data[3] .power_up = "low";

dffeas \data[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_2),
	.prn(vcc));
defparam \data[2] .is_wysiwyg = "true";
defparam \data[2] .power_up = "low";

dffeas \data[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_1),
	.prn(vcc));
defparam \data[1] .is_wysiwyg = "true";
defparam \data[1] .power_up = "low";

dffeas \data[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_0),
	.prn(vcc));
defparam \data[0] .is_wysiwyg = "true";
defparam \data[0] .power_up = "low";

dffeas \data[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_7),
	.prn(vcc));
defparam \data[7] .is_wysiwyg = "true";
defparam \data[7] .power_up = "low";

dffeas \data[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_6),
	.prn(vcc));
defparam \data[6] .is_wysiwyg = "true";
defparam \data[6] .power_up = "low";

dffeas \data[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_5),
	.prn(vcc));
defparam \data[5] .is_wysiwyg = "true";
defparam \data[5] .power_up = "low";

dffeas \data[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\data~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(data_4),
	.prn(vcc));
defparam \data[4] .is_wysiwyg = "true";
defparam \data[4] .power_up = "low";

dffeas err(
	.clk(mac_rx_clock_connection_clk),
	.d(\err~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(\data[7]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.q(err1),
	.prn(vcc));
defparam err.is_wysiwyg = "true";
defparam err.power_up = "low";

cyclonev_lcell_comb \en~0 (
	.dataa(!\U_LBR|Selector1~0_combout ),
	.datab(!\U_LBR|state.STM_TYPE_FRM_READ~q ),
	.datac(!gm_rx_en_i_reg),
	.datad(!\U_LBR|ff_gmii_reg~q ),
	.datae(!dreg_1),
	.dataf(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datag(!packet_in_progress),
	.cin(gnd),
	.sharein(gnd),
	.combout(\en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \en~0 .extended_lut = "on";
defparam \en~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \en~0 .shared_arith = "off";

cyclonev_lcell_comb \data[7]~0 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_LBR|ff_gmii_reg~q ),
	.datac(!\U_LBR|state.STM_TYPE_FRM_READ~q ),
	.datad(!\U_LBFF|aempty_flag~q ),
	.datae(!\U_LBR|state.STM_TYPE_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data[7]~0 .extended_lut = "off";
defparam \data[7]~0 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \data[7]~0 .shared_arith = "off";

dffeas \data_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[3]~q ),
	.prn(vcc));
defparam \data_reg[3] .is_wysiwyg = "true";
defparam \data_reg[3] .power_up = "low";

cyclonev_lcell_comb \data~1 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!gm_rx_d_i_reg_3),
	.datad(!\data_reg[3]~q ),
	.datae(!mii_rxd_o_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~1 .extended_lut = "off";
defparam \data~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~1 .shared_arith = "off";

dffeas \data_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[2]~q ),
	.prn(vcc));
defparam \data_reg[2] .is_wysiwyg = "true";
defparam \data_reg[2] .power_up = "low";

cyclonev_lcell_comb \data~2 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!gm_rx_d_i_reg_2),
	.datad(!\data_reg[2]~q ),
	.datae(!mii_rxd_o_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~2 .extended_lut = "off";
defparam \data~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~2 .shared_arith = "off";

dffeas \data_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[1]~q ),
	.prn(vcc));
defparam \data_reg[1] .is_wysiwyg = "true";
defparam \data_reg[1] .power_up = "low";

cyclonev_lcell_comb \data~3 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!gm_rx_d_i_reg_1),
	.datad(!\data_reg[1]~q ),
	.datae(!mii_rxd_o_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~3 .extended_lut = "off";
defparam \data~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~3 .shared_arith = "off";

dffeas \data_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[0]~q ),
	.prn(vcc));
defparam \data_reg[0] .is_wysiwyg = "true";
defparam \data_reg[0] .power_up = "low";

cyclonev_lcell_comb \data~4 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!gm_rx_d_i_reg_0),
	.datad(!\data_reg[0]~q ),
	.datae(!mii_rxd_o_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~4 .extended_lut = "off";
defparam \data~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~4 .shared_arith = "off";

dffeas \data_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[7]~q ),
	.prn(vcc));
defparam \data_reg[7] .is_wysiwyg = "true";
defparam \data_reg[7] .power_up = "low";

cyclonev_lcell_comb \data~5 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!\data_reg[7]~q ),
	.datad(!gm_rx_d_i_reg_7),
	.datae(!mii_rxd_o_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~5 .extended_lut = "off";
defparam \data~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~5 .shared_arith = "off";

dffeas \data_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[6]~q ),
	.prn(vcc));
defparam \data_reg[6] .is_wysiwyg = "true";
defparam \data_reg[6] .power_up = "low";

cyclonev_lcell_comb \data~6 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!\data_reg[6]~q ),
	.datad(!gm_rx_d_i_reg_6),
	.datae(!mii_rxd_o_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~6 .extended_lut = "off";
defparam \data~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~6 .shared_arith = "off";

dffeas \data_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[5]~q ),
	.prn(vcc));
defparam \data_reg[5] .is_wysiwyg = "true";
defparam \data_reg[5] .power_up = "low";

cyclonev_lcell_comb \data~7 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!\data_reg[5]~q ),
	.datad(!gm_rx_d_i_reg_5),
	.datae(!mii_rxd_o_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~7 .extended_lut = "off";
defparam \data~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~7 .shared_arith = "off";

dffeas \data_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\data_reg[4]~q ),
	.prn(vcc));
defparam \data_reg[4] .is_wysiwyg = "true";
defparam \data_reg[4] .power_up = "low";

cyclonev_lcell_comb \data~8 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!\data_reg[4]~q ),
	.datad(!gm_rx_d_i_reg_4),
	.datae(!mii_rxd_o_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data~8 .extended_lut = "off";
defparam \data~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \data~8 .shared_arith = "off";

dffeas err_reg(
	.clk(mac_rx_clock_connection_clk),
	.d(\U_LBFF|U_RAM|altsyncram_component|auto_generated|q_b[9] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(!\U_LBFF|aempty_low_det~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\err_reg~q ),
	.prn(vcc));
defparam err_reg.is_wysiwyg = "true";
defparam err_reg.power_up = "low";

cyclonev_lcell_comb \err~0 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!dreg_1),
	.datac(!\err_reg~q ),
	.datad(!gm_rx_err_i_reg),
	.datae(!mii_rxerr_o),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\err~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \err~0 .extended_lut = "off";
defparam \err~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \err~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_21 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_21 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_21 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_a_fifo_24 (
	ff_gmii_reg,
	q_b_8,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_9,
	altera_tse_reset_synchronizer_chain_out,
	altera_tse_reset_synchronizer_chain_out1,
	tx_en_s_1,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	stateSTM_TYPE_FRM_READ,
	aempty_flag1,
	Selector1,
	aempty_low_det1,
	Selector11,
	afull_flag1,
	ff_wren,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	ff_gmii_reg;
output 	q_b_8;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_9;
input 	altera_tse_reset_synchronizer_chain_out;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	tx_en_s_1;
input 	rd_14_4;
input 	rd_14_0;
input 	rd_14_5;
input 	rd_14_1;
input 	rd_14_6;
input 	rd_14_2;
input 	rd_14_7;
input 	rd_14_3;
input 	tx_err;
input 	stateSTM_TYPE_FRM_READ;
output 	aempty_flag1;
input 	Selector1;
output 	aempty_low_det1;
input 	Selector11;
output 	afull_flag1;
input 	ff_wren;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_WRT|b_out[0]~q ;
wire \U_WRT|b_out[1]~q ;
wire \U_WRT|b_out[2]~q ;
wire \U_WRT|b_out[3]~q ;
wire \U_WRT|b_out[4]~q ;
wire \U_RD|b_out[0]~q ;
wire \U_RD|b_out[1]~q ;
wire \U_RD|b_out[2]~q ;
wire \U_RD|b_out[3]~q ;
wire \U_RD|b_out[4]~q ;
wire \U_SYNC_WR_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ;
wire \U_WRT|g_out[0]~q ;
wire \U_WRT|g_out[1]~q ;
wire \U_WRT|g_out[2]~q ;
wire \U_WRT|g_out[3]~q ;
wire \U_WRT|g_out[4]~q ;
wire \U_SYNC_RD_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_RD_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_RD_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_RD_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_RD_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ;
wire \U_RD|g_out[4]~q ;
wire \U_RD|g_out[3]~q ;
wire \U_RD|g_out[2]~q ;
wire \U_RD|g_out[1]~q ;
wire \U_RD|g_out[0]~q ;
wire \ff_wr_binval[0]~combout ;
wire \wr_b_rptr[0]~q ;
wire \ptr_rck_diff[0]~1_sumout ;
wire \ff_wr_binval[0]~0_combout ;
wire \wr_b_rptr[1]~q ;
wire \ptr_rck_diff[0]~2 ;
wire \ptr_rck_diff[0]~3 ;
wire \ptr_rck_diff[1]~5_sumout ;
wire \ff_wr_binval[1]~1_combout ;
wire \wr_b_rptr[2]~q ;
wire \ptr_rck_diff[1]~6 ;
wire \ptr_rck_diff[1]~7 ;
wire \ptr_rck_diff[2]~9_sumout ;
wire \ff_wr_binval[3]~2_combout ;
wire \wr_b_rptr[3]~q ;
wire \ptr_rck_diff[2]~10 ;
wire \ptr_rck_diff[2]~11 ;
wire \ptr_rck_diff[3]~13_sumout ;
wire \wr_b_rptr[4]~q ;
wire \ptr_rck_diff[3]~14 ;
wire \ptr_rck_diff[3]~15 ;
wire \ptr_rck_diff[4]~17_sumout ;
wire \LessThan1~0_combout ;
wire \aempty_low_det~0_combout ;
wire \rd_b_wptr[4]~q ;
wire \ff_rd_binval[3]~0_combout ;
wire \rd_b_wptr[3]~q ;
wire \ff_rd_binval[1]~1_combout ;
wire \rd_b_wptr[2]~q ;
wire \ff_rd_binval[0]~2_combout ;
wire \rd_b_wptr[1]~q ;
wire \ff_rd_binval[0]~combout ;
wire \rd_b_wptr[0]~q ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~1_sumout ;
wire \ptr_wck_diff[4]~q ;
wire \Add0~5_sumout ;
wire \ptr_wck_diff[3]~q ;
wire \Add0~9_sumout ;
wire \ptr_wck_diff[2]~q ;
wire \Add0~13_sumout ;
wire \ptr_wck_diff[1]~q ;
wire \Add0~17_sumout ;
wire \ptr_wck_diff[0]~q ;
wire \LessThan0~0_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_1 U_SYNC_WR_G_PTR(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_0(\U_SYNC_WR_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_01(\U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_02(\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_03(\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_04(\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle U_SYNC_RD_G_PTR(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(\U_SYNC_RD_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_01(\U_SYNC_RD_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_02(\U_SYNC_RD_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_03(\U_SYNC_RD_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_04(\U_SYNC_RD_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ),
	.g_out_4(\U_RD|g_out[4]~q ),
	.g_out_3(\U_RD|g_out[3]~q ),
	.g_out_2(\U_RD|g_out[2]~q ),
	.g_out_1(\U_RD|g_out[1]~q ),
	.g_out_0(\U_RD|g_out[0]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt U_RD(
	.ff_gmii_reg(ff_gmii_reg),
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.stateSTM_TYPE_FRM_READ(stateSTM_TYPE_FRM_READ),
	.Selector1(Selector1),
	.Selector11(Selector11),
	.b_out_0(\U_RD|b_out[0]~q ),
	.b_out_1(\U_RD|b_out[1]~q ),
	.b_out_2(\U_RD|b_out[2]~q ),
	.b_out_3(\U_RD|b_out[3]~q ),
	.b_out_4(\U_RD|b_out[4]~q ),
	.g_out_4(\U_RD|g_out[4]~q ),
	.g_out_3(\U_RD|g_out[3]~q ),
	.g_out_2(\U_RD|g_out[2]~q ),
	.g_out_1(\U_RD|g_out[1]~q ),
	.g_out_0(\U_RD|g_out[0]~q ),
	.clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_1 U_WRT(
	.reset(altera_tse_reset_synchronizer_chain_out),
	.ff_wren(ff_wren),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_sdpm_altsyncram U_RAM(
	.q_b_8(q_b_8),
	.q_b_3(q_b_3),
	.q_b_2(q_b_2),
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.q_b_7(q_b_7),
	.q_b_6(q_b_6),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_9(q_b_9),
	.tx_en_s_1(tx_en_s_1),
	.rd_14_4(rd_14_4),
	.rd_14_0(rd_14_0),
	.rd_14_5(rd_14_5),
	.rd_14_1(rd_14_1),
	.rd_14_6(rd_14_6),
	.rd_14_2(rd_14_2),
	.rd_14_7(rd_14_7),
	.rd_14_3(rd_14_3),
	.tx_err(tx_err),
	.ff_wren(ff_wren),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_01(\U_RD|b_out[0]~q ),
	.b_out_11(\U_RD|b_out[1]~q ),
	.b_out_21(\U_RD|b_out[2]~q ),
	.b_out_31(\U_RD|b_out[3]~q ),
	.b_out_41(\U_RD|b_out[4]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

dffeas aempty_flag(
	.clk(mac_rx_clock_connection_clk),
	.d(\LessThan1~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(aempty_flag1),
	.prn(vcc));
defparam aempty_flag.is_wysiwyg = "true";
defparam aempty_flag.power_up = "low";

dffeas aempty_low_det(
	.clk(mac_rx_clock_connection_clk),
	.d(\aempty_low_det~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(aempty_low_det1),
	.prn(vcc));
defparam aempty_low_det.is_wysiwyg = "true";
defparam aempty_low_det.power_up = "low";

dffeas afull_flag(
	.clk(mac_tx_clock_connection_clk),
	.d(\LessThan0~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(afull_flag1),
	.prn(vcc));
defparam afull_flag.is_wysiwyg = "true";
defparam afull_flag.power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0] (
	.dataa(!\U_SYNC_WR_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datad(!\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.datae(!\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0] .extended_lut = "off";
defparam \ff_wr_binval[0] .lut_mask = 64'h9669699696696996;
defparam \ff_wr_binval[0] .shared_arith = "off";

dffeas \wr_b_rptr[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_wr_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[0]~q ),
	.prn(vcc));
defparam \wr_b_rptr[0] .is_wysiwyg = "true";
defparam \wr_b_rptr[0] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[0]~q ),
	.datad(!\U_RD|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\ptr_rck_diff[0]~1_sumout ),
	.cout(\ptr_rck_diff[0]~2 ),
	.shareout(\ptr_rck_diff[0]~3 ));
defparam \ptr_rck_diff[0]~1 .extended_lut = "off";
defparam \ptr_rck_diff[0]~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[0]~1 .shared_arith = "on";

cyclonev_lcell_comb \ff_wr_binval[0]~0 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.datad(!\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0]~0 .extended_lut = "off";
defparam \ff_wr_binval[0]~0 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[0]~0 .shared_arith = "off";

dffeas \wr_b_rptr[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_wr_binval[0]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[1]~q ),
	.prn(vcc));
defparam \wr_b_rptr[1] .is_wysiwyg = "true";
defparam \wr_b_rptr[1] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[1]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[1]~q ),
	.datad(!\U_RD|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[0]~2 ),
	.sharein(\ptr_rck_diff[0]~3 ),
	.combout(),
	.sumout(\ptr_rck_diff[1]~5_sumout ),
	.cout(\ptr_rck_diff[1]~6 ),
	.shareout(\ptr_rck_diff[1]~7 ));
defparam \ptr_rck_diff[1]~5 .extended_lut = "off";
defparam \ptr_rck_diff[1]~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[1]~5 .shared_arith = "on";

cyclonev_lcell_comb \ff_wr_binval[1]~1 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[1]~1 .extended_lut = "off";
defparam \ff_wr_binval[1]~1 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[1]~1 .shared_arith = "off";

dffeas \wr_b_rptr[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_wr_binval[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[2]~q ),
	.prn(vcc));
defparam \wr_b_rptr[2] .is_wysiwyg = "true";
defparam \wr_b_rptr[2] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[2]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[2]~q ),
	.datad(!\U_RD|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[1]~6 ),
	.sharein(\ptr_rck_diff[1]~7 ),
	.combout(),
	.sumout(\ptr_rck_diff[2]~9_sumout ),
	.cout(\ptr_rck_diff[2]~10 ),
	.shareout(\ptr_rck_diff[2]~11 ));
defparam \ptr_rck_diff[2]~9 .extended_lut = "off";
defparam \ptr_rck_diff[2]~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[2]~9 .shared_arith = "on";

cyclonev_lcell_comb \ff_wr_binval[3]~2 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~2 .extended_lut = "off";
defparam \ff_wr_binval[3]~2 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[3]~2 .shared_arith = "off";

dffeas \wr_b_rptr[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_wr_binval[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[3]~q ),
	.prn(vcc));
defparam \wr_b_rptr[3] .is_wysiwyg = "true";
defparam \wr_b_rptr[3] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[3]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[3]~q ),
	.datad(!\U_RD|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[2]~10 ),
	.sharein(\ptr_rck_diff[2]~11 ),
	.combout(),
	.sumout(\ptr_rck_diff[3]~13_sumout ),
	.cout(\ptr_rck_diff[3]~14 ),
	.shareout(\ptr_rck_diff[3]~15 ));
defparam \ptr_rck_diff[3]~13 .extended_lut = "off";
defparam \ptr_rck_diff[3]~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[3]~13 .shared_arith = "on";

dffeas \wr_b_rptr[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[4]~q ),
	.prn(vcc));
defparam \wr_b_rptr[4] .is_wysiwyg = "true";
defparam \wr_b_rptr[4] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[4]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[4]~q ),
	.datad(!\U_RD|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[3]~14 ),
	.sharein(\ptr_rck_diff[3]~15 ),
	.combout(),
	.sumout(\ptr_rck_diff[4]~17_sumout ),
	.cout(),
	.shareout());
defparam \ptr_rck_diff[4]~17 .extended_lut = "off";
defparam \ptr_rck_diff[4]~17 .lut_mask = 64'h0000000000000FF0;
defparam \ptr_rck_diff[4]~17 .shared_arith = "on";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!\ptr_rck_diff[0]~1_sumout ),
	.datab(!\ptr_rck_diff[1]~5_sumout ),
	.datac(!\ptr_rck_diff[2]~9_sumout ),
	.datad(!\ptr_rck_diff[3]~13_sumout ),
	.datae(!\ptr_rck_diff[4]~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \aempty_low_det~0 (
	.dataa(!aempty_flag1),
	.datab(!aempty_low_det1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_low_det~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_low_det~0 .extended_lut = "off";
defparam \aempty_low_det~0 .lut_mask = 64'h7777777777777777;
defparam \aempty_low_det~0 .shared_arith = "off";

dffeas \rd_b_wptr[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_SYNC_RD_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[4]~q ),
	.prn(vcc));
defparam \rd_b_wptr[4] .is_wysiwyg = "true";
defparam \rd_b_wptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[3]~0 (
	.dataa(!\U_SYNC_RD_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_RD_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[3]~0 .extended_lut = "off";
defparam \ff_rd_binval[3]~0 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[3]~0 .shared_arith = "off";

dffeas \rd_b_wptr[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_rd_binval[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[3]~q ),
	.prn(vcc));
defparam \rd_b_wptr[3] .is_wysiwyg = "true";
defparam \rd_b_wptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[1]~1 (
	.dataa(!\ff_rd_binval[3]~0_combout ),
	.datab(!\U_SYNC_RD_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[1]~1 .extended_lut = "off";
defparam \ff_rd_binval[1]~1 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[1]~1 .shared_arith = "off";

dffeas \rd_b_wptr[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_rd_binval[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[2]~q ),
	.prn(vcc));
defparam \rd_b_wptr[2] .is_wysiwyg = "true";
defparam \rd_b_wptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[0]~2 (
	.dataa(!\ff_rd_binval[1]~1_combout ),
	.datab(!\U_SYNC_RD_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[0]~2 .extended_lut = "off";
defparam \ff_rd_binval[0]~2 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[0]~2 .shared_arith = "off";

dffeas \rd_b_wptr[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_rd_binval[0]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[1]~q ),
	.prn(vcc));
defparam \rd_b_wptr[1] .is_wysiwyg = "true";
defparam \rd_b_wptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[0] (
	.dataa(!\ff_rd_binval[0]~2_combout ),
	.datab(!\U_SYNC_RD_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[0] .extended_lut = "off";
defparam \ff_rd_binval[0] .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[0] .shared_arith = "off";

dffeas \rd_b_wptr[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_rd_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[0]~q ),
	.prn(vcc));
defparam \rd_b_wptr[0] .is_wysiwyg = "true";
defparam \rd_b_wptr[0] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[0]~q ),
	.datad(!\U_WRT|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[1]~q ),
	.datad(!\U_WRT|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[2]~q ),
	.datad(!\U_WRT|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[3]~q ),
	.datad(!\U_WRT|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[4]~q ),
	.datad(!\U_WRT|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000000000000FF0;
defparam \Add0~1 .shared_arith = "on";

dffeas \ptr_wck_diff[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[4]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[4] .is_wysiwyg = "true";
defparam \ptr_wck_diff[4] .power_up = "low";

dffeas \ptr_wck_diff[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[3]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[3] .is_wysiwyg = "true";
defparam \ptr_wck_diff[3] .power_up = "low";

dffeas \ptr_wck_diff[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[2]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[2] .is_wysiwyg = "true";
defparam \ptr_wck_diff[2] .power_up = "low";

dffeas \ptr_wck_diff[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[1]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[1] .is_wysiwyg = "true";
defparam \ptr_wck_diff[1] .power_up = "low";

dffeas \ptr_wck_diff[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[0]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[0] .is_wysiwyg = "true";
defparam \ptr_wck_diff[0] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\ptr_wck_diff[4]~q ),
	.datab(!\ptr_wck_diff[3]~q ),
	.datac(!\ptr_wck_diff[2]~q ),
	.datad(!\ptr_wck_diff[1]~q ),
	.datae(!\ptr_wck_diff[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan0~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	dreg_01,
	dreg_02,
	dreg_03,
	dreg_04,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
output 	dreg_01;
output 	dreg_02;
output 	dreg_03;
output 	dreg_04;
input 	g_out_4;
input 	g_out_3;
input 	g_out_2;
input 	g_out_1;
input 	g_out_0;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_26 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.g_out_4(g_out_4),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_25 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_01),
	.g_out_3(g_out_3),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_24 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_02),
	.g_out_2(g_out_2),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_23 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_03),
	.g_out_1(g_out_1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_22 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_04),
	.g_out_0(g_out_0),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_22 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_0,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_0;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_22 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_0),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_22 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_23 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_23 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_23 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_24 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_2,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_2;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_24 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_2),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_24 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_25 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_3,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_3;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_25 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_3),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_25 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_26 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_4,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_4;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_26 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_4),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_26 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_1 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	dreg_01,
	dreg_02,
	dreg_03,
	dreg_04,
	g_out_0,
	g_out_1,
	g_out_2,
	g_out_3,
	g_out_4,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
output 	dreg_01;
output 	dreg_02;
output 	dreg_03;
output 	dreg_04;
input 	g_out_0;
input 	g_out_1;
input 	g_out_2;
input 	g_out_3;
input 	g_out_4;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_31 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_04),
	.g_out_4(g_out_4),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_30 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_03),
	.g_out_3(g_out_3),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_29 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_02),
	.g_out_2(g_out_2),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_28 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_01),
	.g_out_1(g_out_1),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_27 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.g_out_0(g_out_0),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_27 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_0,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_0;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_27 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_0),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_27 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_28 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_28 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_28 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_29 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_2,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_2;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_29 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_2),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_29 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_30 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_3,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_3;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_30 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_3),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_30 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_31 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	g_out_4,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	g_out_4;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_31 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(g_out_4),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_31 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt (
	ff_gmii_reg,
	reset,
	stateSTM_TYPE_FRM_READ,
	Selector1,
	Selector11,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	ff_gmii_reg;
input 	reset;
input 	stateSTM_TYPE_FRM_READ;
input 	Selector1;
input 	Selector11;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	g_out_4;
output 	g_out_3;
output 	g_out_2;
output 	g_out_1;
output 	g_out_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \b_int[0]~4_combout ;
wire \b_int[0]~q ;
wire \b_out[0]~0_combout ;
wire \Add0~0_combout ;
wire \b_int[1]~q ;
wire \b_int[2]~0_combout ;
wire \b_int[2]~1_combout ;
wire \b_int[2]~q ;
wire \b_int[3]~2_combout ;
wire \b_int[3]~q ;
wire \b_int[4]~3_combout ;
wire \b_int[4]~q ;
wire \gry_grayval[3]~combout ;
wire \gry_grayval[2]~combout ;
wire \gry_grayval[1]~combout ;


dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \g_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[3] (
	.clk(clk),
	.d(\gry_grayval[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[2] (
	.clk(clk),
	.d(\gry_grayval[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[1] (
	.clk(clk),
	.d(\gry_grayval[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[0] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

cyclonev_lcell_comb \b_int[0]~4 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[0]~4 .extended_lut = "off";
defparam \b_int[0]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_int[0]~4 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6666666666666666;
defparam \Add0~0 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(Selector11),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \b_int[2]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[2]~0 .extended_lut = "off";
defparam \b_int[2]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \b_int[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \b_int[2]~1 (
	.dataa(!ff_gmii_reg),
	.datab(!stateSTM_TYPE_FRM_READ),
	.datac(!Selector1),
	.datad(!\b_int[2]~q ),
	.datae(!\b_int[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[2]~1 .extended_lut = "off";
defparam \b_int[2]~1 .lut_mask = 64'h9669699696696996;
defparam \b_int[2]~1 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\b_int[2]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

cyclonev_lcell_comb \b_int[3]~2 (
	.dataa(!ff_gmii_reg),
	.datab(!stateSTM_TYPE_FRM_READ),
	.datac(!Selector1),
	.datad(!\b_int[2]~q ),
	.datae(!\b_int[3]~q ),
	.dataf(!\b_int[2]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[3]~2 .extended_lut = "off";
defparam \b_int[3]~2 .lut_mask = 64'h6996966996696996;
defparam \b_int[3]~2 .shared_arith = "off";

dffeas \b_int[3] (
	.clk(clk),
	.d(\b_int[3]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \b_int[4]~3 (
	.dataa(!Selector11),
	.datab(!\b_int[2]~q ),
	.datac(!\b_int[3]~q ),
	.datad(!\b_int[4]~q ),
	.datae(!\b_int[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[4]~3 .extended_lut = "off";
defparam \b_int[4]~3 .lut_mask = 64'h9669699696696996;
defparam \b_int[4]~3 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\b_int[4]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \gry_grayval[3] (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[3] .extended_lut = "off";
defparam \gry_grayval[3] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[3] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[2] (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[2] .extended_lut = "off";
defparam \gry_grayval[2] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[2] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[1] (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[1] .extended_lut = "off";
defparam \gry_grayval[1] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[1] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_1 (
	reset,
	ff_wren,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	g_out_0,
	g_out_1,
	g_out_2,
	g_out_3,
	g_out_4,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	ff_wren;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	g_out_0;
output 	g_out_1;
output 	g_out_2;
output 	g_out_3;
output 	g_out_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \b_int[0]~3_combout ;
wire \b_int[0]~q ;
wire \b_out[0]~0_combout ;
wire \Add0~0_combout ;
wire \b_int[1]~q ;
wire \b_int[2]~0_combout ;
wire \b_int[2]~q ;
wire \b_int[3]~1_combout ;
wire \b_int[3]~q ;
wire \b_int[4]~2_combout ;
wire \b_int[4]~q ;
wire \gry_grayval[1]~combout ;
wire \gry_grayval[2]~combout ;
wire \gry_grayval[3]~combout ;


dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \g_out[0] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

dffeas \g_out[1] (
	.clk(clk),
	.d(\gry_grayval[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[2] (
	.clk(clk),
	.d(\gry_grayval[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[3] (
	.clk(clk),
	.d(\gry_grayval[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

cyclonev_lcell_comb \b_int[0]~3 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[0]~3 .extended_lut = "off";
defparam \b_int[0]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_int[0]~3 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int[0]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h6666666666666666;
defparam \Add0~0 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ff_wren),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \b_int[2]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(!\b_int[2]~q ),
	.datad(!ff_wren),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[2]~0 .extended_lut = "off";
defparam \b_int[2]~0 .lut_mask = 64'h6996699669966996;
defparam \b_int[2]~0 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\b_int[2]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

cyclonev_lcell_comb \b_int[3]~1 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(!\b_int[2]~q ),
	.datad(!\b_int[3]~q ),
	.datae(!ff_wren),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[3]~1 .extended_lut = "off";
defparam \b_int[3]~1 .lut_mask = 64'h9669699696696996;
defparam \b_int[3]~1 .shared_arith = "off";

dffeas \b_int[3] (
	.clk(clk),
	.d(\b_int[3]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \b_int[4]~2 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(!\b_int[2]~q ),
	.datad(!\b_int[3]~q ),
	.datae(!\b_int[4]~q ),
	.dataf(!ff_wren),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int[4]~2 .extended_lut = "off";
defparam \b_int[4]~2 .lut_mask = 64'h6996966996696996;
defparam \b_int[4]~2 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\b_int[4]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \gry_grayval[1] (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[1] .extended_lut = "off";
defparam \gry_grayval[1] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[1] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[2] (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[2] .extended_lut = "off";
defparam \gry_grayval[2] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[2] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[3] (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[3] .extended_lut = "off";
defparam \gry_grayval[3] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[3] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_sdpm_altsyncram (
	q_b_8,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_0,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_9,
	tx_en_s_1,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	ff_wren,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_01,
	b_out_11,
	b_out_21,
	b_out_31,
	b_out_41,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_8;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
output 	q_b_0;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_9;
input 	tx_en_s_1;
input 	rd_14_4;
input 	rd_14_0;
input 	rd_14_5;
input 	rd_14_1;
input 	rd_14_6;
input 	rd_14_2;
input 	rd_14_7;
input 	rd_14_3;
input 	tx_err;
input 	ff_wren;
input 	b_out_0;
input 	b_out_1;
input 	b_out_2;
input 	b_out_3;
input 	b_out_4;
input 	b_out_01;
input 	b_out_11;
input 	b_out_21;
input 	b_out_31;
input 	b_out_41;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_1 altsyncram_component(
	.q_b({q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_unconnected_wire_35,q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,
q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,
q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,tx_err,tx_en_s_1,rd_14_7,rd_14_6,rd_14_5,rd_14_4,rd_14_3,rd_14_2,rd_14_1,rd_14_0}),
	.wren_a(ff_wren),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,b_out_4,b_out_3,b_out_2,b_out_1,b_out_0}),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,b_out_41,b_out_31,b_out_21,b_out_11,b_out_01}),
	.clock0(mac_tx_clock_connection_clk),
	.clock1(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altsyncram_1 (
	q_b,
	data_a,
	wren_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	[39:0] data_a;
input 	wren_a;
input 	[10:0] address_a;
input 	[10:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_2vl1 auto_generated(
	.q_b({q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0),
	.clock1(clock1));

endmodule

module IoTOctopus_QSYS_altsyncram_2vl1 (
	q_b,
	data_a,
	wren_a,
	address_a,
	address_b,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[9:0] q_b;
input 	[9:0] data_a;
input 	wren_a;
input 	[4:0] address_a;
input 	[4:0] address_b;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 10;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 10;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 10;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 10;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 10;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 10;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 10;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 10;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 10;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_loopback_ff:U_LBFF|altera_tse_a_fifo_24:U_LBFF|altera_tse_sdpm_altsyncram:U_RAM|altsyncram:altsyncram_component|altsyncram_2vl1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 10;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

endmodule

module IoTOctopus_QSYS_altera_tse_lb_read_cntl (
	ff_gmii_reg1,
	ff_gmii_en,
	reset,
	stateSTM_TYPE_FRM_READ,
	aempty_flag,
	stateSTM_TYPE_IDLE,
	Selector1,
	aempty_low_det,
	Selector11,
	clk)/* synthesis synthesis_greybox=1 */;
output 	ff_gmii_reg1;
input 	ff_gmii_en;
input 	reset;
output 	stateSTM_TYPE_FRM_READ;
input 	aempty_flag;
output 	stateSTM_TYPE_IDLE;
output 	Selector1;
input 	aempty_low_det;
output 	Selector11;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nextstate.STM_TYPE_NEXT_FRM~0_combout ;
wire \state.STM_TYPE_NEXT_FRM~q ;
wire \Selector0~0_combout ;


dffeas ff_gmii_reg(
	.clk(clk),
	.d(ff_gmii_en),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(!aempty_low_det),
	.sload(gnd),
	.ena(vcc),
	.q(ff_gmii_reg1),
	.prn(vcc));
defparam ff_gmii_reg.is_wysiwyg = "true";
defparam ff_gmii_reg.power_up = "low";

dffeas \state.STM_TYPE_FRM_READ (
	.clk(clk),
	.d(Selector11),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateSTM_TYPE_FRM_READ),
	.prn(vcc));
defparam \state.STM_TYPE_FRM_READ .is_wysiwyg = "true";
defparam \state.STM_TYPE_FRM_READ .power_up = "low";

dffeas \state.STM_TYPE_IDLE (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateSTM_TYPE_IDLE),
	.prn(vcc));
defparam \state.STM_TYPE_IDLE .is_wysiwyg = "true";
defparam \state.STM_TYPE_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!aempty_flag),
	.datab(!stateSTM_TYPE_IDLE),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!ff_gmii_reg1),
	.datab(!stateSTM_TYPE_FRM_READ),
	.datac(!aempty_flag),
	.datad(!stateSTM_TYPE_IDLE),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \nextstate.STM_TYPE_NEXT_FRM~0 (
	.dataa(!ff_gmii_reg1),
	.datab(!stateSTM_TYPE_FRM_READ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nextstate.STM_TYPE_NEXT_FRM~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nextstate.STM_TYPE_NEXT_FRM~0 .extended_lut = "off";
defparam \nextstate.STM_TYPE_NEXT_FRM~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nextstate.STM_TYPE_NEXT_FRM~0 .shared_arith = "off";

dffeas \state.STM_TYPE_NEXT_FRM (
	.clk(clk),
	.d(\nextstate.STM_TYPE_NEXT_FRM~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYPE_NEXT_FRM~q ),
	.prn(vcc));
defparam \state.STM_TYPE_NEXT_FRM .is_wysiwyg = "true";
defparam \state.STM_TYPE_NEXT_FRM .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!aempty_flag),
	.datab(!stateSTM_TYPE_IDLE),
	.datac(!\state.STM_TYPE_NEXT_FRM~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Selector0~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_lb_wrt_cntl (
	altera_tse_reset_synchronizer_chain_out,
	tx_en_s_1,
	afull_flag,
	ff_wren,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
input 	tx_en_s_1;
input 	afull_flag;
output 	ff_wren;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_LOOPBACK_ENA|std_sync_no_cut|dreg[1]~q ;
wire \nextstate.STM_TYPE_NEXT_FRM~0_combout ;
wire \state.STM_TYPE_NEXT_FRM~q ;
wire \Selector0~0_combout ;
wire \state.STM_TYPE_IDLE~q ;
wire \Selector1~0_combout ;
wire \state.STM_TYPE_LOOP_ENA~q ;
wire \Selector2~0_combout ;
wire \state.STM_TYPE_FRM_WRT~q ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_32 U_SYNC_LOOPBACK_ENA(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_LOOPBACK_ENA|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

cyclonev_lcell_comb \ff_wren~0 (
	.dataa(!tx_en_s_1),
	.datab(!\state.STM_TYPE_FRM_WRT~q ),
	.datac(!\state.STM_TYPE_NEXT_FRM~q ),
	.datad(!afull_flag),
	.datae(!\state.STM_TYPE_LOOP_ENA~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_wren),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wren~0 .extended_lut = "off";
defparam \ff_wren~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \ff_wren~0 .shared_arith = "off";

cyclonev_lcell_comb \nextstate.STM_TYPE_NEXT_FRM~0 (
	.dataa(!tx_en_s_1),
	.datab(!\state.STM_TYPE_FRM_WRT~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nextstate.STM_TYPE_NEXT_FRM~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nextstate.STM_TYPE_NEXT_FRM~0 .extended_lut = "off";
defparam \nextstate.STM_TYPE_NEXT_FRM~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nextstate.STM_TYPE_NEXT_FRM~0 .shared_arith = "off";

dffeas \state.STM_TYPE_NEXT_FRM (
	.clk(mac_tx_clock_connection_clk),
	.d(\nextstate.STM_TYPE_NEXT_FRM~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYPE_NEXT_FRM~q ),
	.prn(vcc));
defparam \state.STM_TYPE_NEXT_FRM .is_wysiwyg = "true";
defparam \state.STM_TYPE_NEXT_FRM .power_up = "low";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!tx_en_s_1),
	.datab(!\state.STM_TYPE_NEXT_FRM~q ),
	.datac(!afull_flag),
	.datad(!\state.STM_TYPE_LOOP_ENA~q ),
	.datae(!\U_SYNC_LOOPBACK_ENA|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\state.STM_TYPE_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hFFD8FFFFFFFFFFFF;
defparam \Selector0~0 .shared_arith = "off";

dffeas \state.STM_TYPE_IDLE (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYPE_IDLE~q ),
	.prn(vcc));
defparam \state.STM_TYPE_IDLE .is_wysiwyg = "true";
defparam \state.STM_TYPE_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!tx_en_s_1),
	.datab(!afull_flag),
	.datac(!\state.STM_TYPE_LOOP_ENA~q ),
	.datad(!\U_SYNC_LOOPBACK_ENA|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYPE_IDLE~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hFFFFBFFFFFFFBFFF;
defparam \Selector1~0 .shared_arith = "off";

dffeas \state.STM_TYPE_LOOP_ENA (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector1~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYPE_LOOP_ENA~q ),
	.prn(vcc));
defparam \state.STM_TYPE_LOOP_ENA .is_wysiwyg = "true";
defparam \state.STM_TYPE_LOOP_ENA .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!tx_en_s_1),
	.datab(!\state.STM_TYPE_FRM_WRT~q ),
	.datac(!afull_flag),
	.datad(!\state.STM_TYPE_LOOP_ENA~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \Selector2~0 .shared_arith = "off";

dffeas \state.STM_TYPE_FRM_WRT (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYPE_FRM_WRT~q ),
	.prn(vcc));
defparam \state.STM_TYPE_FRM_WRT .is_wysiwyg = "true";
defparam \state.STM_TYPE_FRM_WRT .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_32 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_32 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_32 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_mii_rx_if (
	mii_rxd_o_3,
	mii_rxd_o_2,
	mii_rxd_o_1,
	mii_rxd_o_0,
	mii_rxd_o_7,
	mii_rxd_o_6,
	mii_rxd_o_5,
	mii_rxd_o_4,
	mii_rxerr_o1,
	reset,
	mii_clk_ena1,
	gm_rx_en_i_reg,
	packet_in_progress1,
	gm_rx_d_i_reg_3,
	gm_rx_d_i_reg_2,
	gm_rx_d_i_reg_1,
	gm_rx_d_i_reg_0,
	gm_rx_err_i_reg,
	rx_clk)/* synthesis synthesis_greybox=1 */;
output 	mii_rxd_o_3;
output 	mii_rxd_o_2;
output 	mii_rxd_o_1;
output 	mii_rxd_o_0;
output 	mii_rxd_o_7;
output 	mii_rxd_o_6;
output 	mii_rxd_o_5;
output 	mii_rxd_o_4;
output 	mii_rxerr_o1;
input 	reset;
output 	mii_clk_ena1;
input 	gm_rx_en_i_reg;
output 	packet_in_progress1;
input 	gm_rx_d_i_reg_3;
input 	gm_rx_d_i_reg_2;
input 	gm_rx_d_i_reg_1;
input 	gm_rx_d_i_reg_0;
input 	gm_rx_err_i_reg;
input 	rx_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mii_rxdv_reg_1~q ;
wire \mii_rxdv_reg_2~q ;
wire \mii_rxd_reg_1[3]~q ;
wire \mii_rxd_reg_1[2]~q ;
wire \mii_rxd_reg_1[1]~q ;
wire \mii_rxd_reg_1[0]~q ;
wire \always2~0_combout ;
wire \always2~1_combout ;
wire \align_pipeline_1_2~0_combout ;
wire \align_pipeline_1_2~q ;
wire \mii_rxd_reg_2[3]~q ;
wire \mii_rxd_o~0_combout ;
wire \mii_rxerr_o~1_combout ;
wire \mii_rxd_reg_2[2]~q ;
wire \mii_rxd_o~1_combout ;
wire \mii_rxd_reg_2[1]~q ;
wire \mii_rxd_o~2_combout ;
wire \mii_rxd_reg_2[0]~q ;
wire \mii_rxd_o~3_combout ;
wire \mii_rxd_o~4_combout ;
wire \mii_rxd_o~5_combout ;
wire \mii_rxd_o~6_combout ;
wire \mii_rxd_o~7_combout ;
wire \mii_rxerr_reg_1~q ;
wire \mii_rxerr_reg_2~q ;
wire \mii_rxerr_o~0_combout ;
wire \mii_clk_ena~0_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~1_combout ;


dffeas \mii_rxd_o[3] (
	.clk(rx_clk),
	.d(\mii_rxd_o~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_3),
	.prn(vcc));
defparam \mii_rxd_o[3] .is_wysiwyg = "true";
defparam \mii_rxd_o[3] .power_up = "low";

dffeas \mii_rxd_o[2] (
	.clk(rx_clk),
	.d(\mii_rxd_o~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_2),
	.prn(vcc));
defparam \mii_rxd_o[2] .is_wysiwyg = "true";
defparam \mii_rxd_o[2] .power_up = "low";

dffeas \mii_rxd_o[1] (
	.clk(rx_clk),
	.d(\mii_rxd_o~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_1),
	.prn(vcc));
defparam \mii_rxd_o[1] .is_wysiwyg = "true";
defparam \mii_rxd_o[1] .power_up = "low";

dffeas \mii_rxd_o[0] (
	.clk(rx_clk),
	.d(\mii_rxd_o~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_0),
	.prn(vcc));
defparam \mii_rxd_o[0] .is_wysiwyg = "true";
defparam \mii_rxd_o[0] .power_up = "low";

dffeas \mii_rxd_o[7] (
	.clk(rx_clk),
	.d(\mii_rxd_o~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_7),
	.prn(vcc));
defparam \mii_rxd_o[7] .is_wysiwyg = "true";
defparam \mii_rxd_o[7] .power_up = "low";

dffeas \mii_rxd_o[6] (
	.clk(rx_clk),
	.d(\mii_rxd_o~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_6),
	.prn(vcc));
defparam \mii_rxd_o[6] .is_wysiwyg = "true";
defparam \mii_rxd_o[6] .power_up = "low";

dffeas \mii_rxd_o[5] (
	.clk(rx_clk),
	.d(\mii_rxd_o~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_5),
	.prn(vcc));
defparam \mii_rxd_o[5] .is_wysiwyg = "true";
defparam \mii_rxd_o[5] .power_up = "low";

dffeas \mii_rxd_o[4] (
	.clk(rx_clk),
	.d(\mii_rxd_o~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxd_o_4),
	.prn(vcc));
defparam \mii_rxd_o[4] .is_wysiwyg = "true";
defparam \mii_rxd_o[4] .power_up = "low";

dffeas mii_rxerr_o(
	.clk(rx_clk),
	.d(\mii_rxerr_o~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\mii_rxerr_o~1_combout ),
	.sload(gnd),
	.ena(mii_clk_ena1),
	.q(mii_rxerr_o1),
	.prn(vcc));
defparam mii_rxerr_o.is_wysiwyg = "true";
defparam mii_rxerr_o.power_up = "low";

dffeas mii_clk_ena(
	.clk(rx_clk),
	.d(\mii_clk_ena~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_clk_ena1),
	.prn(vcc));
defparam mii_clk_ena.is_wysiwyg = "true";
defparam mii_clk_ena.power_up = "low";

dffeas packet_in_progress(
	.clk(rx_clk),
	.d(\packet_in_progress~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(packet_in_progress1),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

dffeas mii_rxdv_reg_1(
	.clk(rx_clk),
	.d(gm_rx_en_i_reg),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxdv_reg_1~q ),
	.prn(vcc));
defparam mii_rxdv_reg_1.is_wysiwyg = "true";
defparam mii_rxdv_reg_1.power_up = "low";

dffeas mii_rxdv_reg_2(
	.clk(rx_clk),
	.d(\mii_rxdv_reg_1~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxdv_reg_2~q ),
	.prn(vcc));
defparam mii_rxdv_reg_2.is_wysiwyg = "true";
defparam mii_rxdv_reg_2.power_up = "low";

dffeas \mii_rxd_reg_1[3] (
	.clk(rx_clk),
	.d(gm_rx_d_i_reg_3),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_1[3]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_1[3] .is_wysiwyg = "true";
defparam \mii_rxd_reg_1[3] .power_up = "low";

dffeas \mii_rxd_reg_1[2] (
	.clk(rx_clk),
	.d(gm_rx_d_i_reg_2),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_1[2]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_1[2] .is_wysiwyg = "true";
defparam \mii_rxd_reg_1[2] .power_up = "low";

dffeas \mii_rxd_reg_1[1] (
	.clk(rx_clk),
	.d(gm_rx_d_i_reg_1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_1[1]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_1[1] .is_wysiwyg = "true";
defparam \mii_rxd_reg_1[1] .power_up = "low";

dffeas \mii_rxd_reg_1[0] (
	.clk(rx_clk),
	.d(gm_rx_d_i_reg_0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_1[0]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_1[0] .is_wysiwyg = "true";
defparam \mii_rxd_reg_1[0] .power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\mii_rxdv_reg_2~q ),
	.datab(!\mii_rxd_reg_1[3]~q ),
	.datac(!\mii_rxd_reg_1[2]~q ),
	.datad(!\mii_rxd_reg_1[1]~q ),
	.datae(!\mii_rxd_reg_1[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \always2~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~1 (
	.dataa(!\mii_rxdv_reg_1~q ),
	.datab(!gm_rx_d_i_reg_3),
	.datac(!gm_rx_d_i_reg_2),
	.datad(!gm_rx_d_i_reg_1),
	.datae(!gm_rx_d_i_reg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \align_pipeline_1_2~0 (
	.dataa(!mii_clk_ena1),
	.datab(!packet_in_progress1),
	.datac(!\align_pipeline_1_2~q ),
	.datad(!\always2~0_combout ),
	.datae(!\always2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\align_pipeline_1_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \align_pipeline_1_2~0 .extended_lut = "off";
defparam \align_pipeline_1_2~0 .lut_mask = 64'hFFFFFF6FFFFFFF6F;
defparam \align_pipeline_1_2~0 .shared_arith = "off";

dffeas align_pipeline_1_2(
	.clk(rx_clk),
	.d(\align_pipeline_1_2~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\align_pipeline_1_2~q ),
	.prn(vcc));
defparam align_pipeline_1_2.is_wysiwyg = "true";
defparam align_pipeline_1_2.power_up = "low";

dffeas \mii_rxd_reg_2[3] (
	.clk(rx_clk),
	.d(\mii_rxd_reg_1[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_2[3]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_2[3] .is_wysiwyg = "true";
defparam \mii_rxd_reg_2[3] .power_up = "low";

cyclonev_lcell_comb \mii_rxd_o~0 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[3]~q ),
	.datad(!\always2~0_combout ),
	.datae(!\mii_rxd_reg_2[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~0 .extended_lut = "off";
defparam \mii_rxd_o~0 .lut_mask = 64'h9F6FFFFF9F6FFFFF;
defparam \mii_rxd_o~0 .shared_arith = "off";

cyclonev_lcell_comb \mii_rxerr_o~1 (
	.dataa(!\mii_rxdv_reg_1~q ),
	.datab(!\always2~1_combout ),
	.datac(!\mii_rxdv_reg_2~q ),
	.datad(!\always2~0_combout ),
	.datae(!\align_pipeline_1_2~q ),
	.dataf(!packet_in_progress1),
	.datag(!gm_rx_en_i_reg),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxerr_o~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxerr_o~1 .extended_lut = "on";
defparam \mii_rxerr_o~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \mii_rxerr_o~1 .shared_arith = "off";

dffeas \mii_rxd_reg_2[2] (
	.clk(rx_clk),
	.d(\mii_rxd_reg_1[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_2[2]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_2[2] .is_wysiwyg = "true";
defparam \mii_rxd_reg_2[2] .power_up = "low";

cyclonev_lcell_comb \mii_rxd_o~1 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[2]~q ),
	.datad(!\always2~0_combout ),
	.datae(!\mii_rxd_reg_2[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~1 .extended_lut = "off";
defparam \mii_rxd_o~1 .lut_mask = 64'h9F6FFFFF9F6FFFFF;
defparam \mii_rxd_o~1 .shared_arith = "off";

dffeas \mii_rxd_reg_2[1] (
	.clk(rx_clk),
	.d(\mii_rxd_reg_1[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_2[1]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_2[1] .is_wysiwyg = "true";
defparam \mii_rxd_reg_2[1] .power_up = "low";

cyclonev_lcell_comb \mii_rxd_o~2 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[1]~q ),
	.datad(!\always2~0_combout ),
	.datae(!\mii_rxd_reg_2[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~2 .extended_lut = "off";
defparam \mii_rxd_o~2 .lut_mask = 64'h9F6FFFFF9F6FFFFF;
defparam \mii_rxd_o~2 .shared_arith = "off";

dffeas \mii_rxd_reg_2[0] (
	.clk(rx_clk),
	.d(\mii_rxd_reg_1[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxd_reg_2[0]~q ),
	.prn(vcc));
defparam \mii_rxd_reg_2[0] .is_wysiwyg = "true";
defparam \mii_rxd_reg_2[0] .power_up = "low";

cyclonev_lcell_comb \mii_rxd_o~3 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[0]~q ),
	.datad(!\always2~0_combout ),
	.datae(!\mii_rxd_reg_2[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~3 .extended_lut = "off";
defparam \mii_rxd_o~3 .lut_mask = 64'h9F6FFFFF9F6FFFFF;
defparam \mii_rxd_o~3 .shared_arith = "off";

cyclonev_lcell_comb \mii_rxd_o~4 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[3]~q ),
	.datad(!gm_rx_d_i_reg_3),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~4 .extended_lut = "off";
defparam \mii_rxd_o~4 .lut_mask = 64'h9FFF6FFF9FFF6FFF;
defparam \mii_rxd_o~4 .shared_arith = "off";

cyclonev_lcell_comb \mii_rxd_o~5 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[2]~q ),
	.datad(!gm_rx_d_i_reg_2),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~5 .extended_lut = "off";
defparam \mii_rxd_o~5 .lut_mask = 64'h9FFF6FFF9FFF6FFF;
defparam \mii_rxd_o~5 .shared_arith = "off";

cyclonev_lcell_comb \mii_rxd_o~6 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[1]~q ),
	.datad(!gm_rx_d_i_reg_1),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~6 .extended_lut = "off";
defparam \mii_rxd_o~6 .lut_mask = 64'h9FFF6FFF9FFF6FFF;
defparam \mii_rxd_o~6 .shared_arith = "off";

cyclonev_lcell_comb \mii_rxd_o~7 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\mii_rxd_reg_1[0]~q ),
	.datad(!gm_rx_d_i_reg_0),
	.datae(!\always2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxd_o~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxd_o~7 .extended_lut = "off";
defparam \mii_rxd_o~7 .lut_mask = 64'h9FFF6FFF9FFF6FFF;
defparam \mii_rxd_o~7 .shared_arith = "off";

dffeas mii_rxerr_reg_1(
	.clk(rx_clk),
	.d(gm_rx_err_i_reg),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxerr_reg_1~q ),
	.prn(vcc));
defparam mii_rxerr_reg_1.is_wysiwyg = "true";
defparam mii_rxerr_reg_1.power_up = "low";

dffeas mii_rxerr_reg_2(
	.clk(rx_clk),
	.d(\mii_rxerr_reg_1~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_rxerr_reg_2~q ),
	.prn(vcc));
defparam mii_rxerr_reg_2.is_wysiwyg = "true";
defparam mii_rxerr_reg_2.power_up = "low";

cyclonev_lcell_comb \mii_rxerr_o~0 (
	.dataa(!packet_in_progress1),
	.datab(!\align_pipeline_1_2~q ),
	.datac(!\always2~0_combout ),
	.datad(!gm_rx_err_i_reg),
	.datae(!\mii_rxerr_reg_1~q ),
	.dataf(!\mii_rxerr_reg_2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_rxerr_o~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_rxerr_o~0 .extended_lut = "off";
defparam \mii_rxerr_o~0 .lut_mask = 64'h96FFFFFFFFFFFFFF;
defparam \mii_rxerr_o~0 .shared_arith = "off";

cyclonev_lcell_comb \mii_clk_ena~0 (
	.dataa(!mii_clk_ena1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_clk_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_clk_ena~0 .extended_lut = "off";
defparam \mii_clk_ena~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \mii_clk_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!gm_rx_en_i_reg),
	.datab(!\mii_rxdv_reg_1~q ),
	.datac(!\align_pipeline_1_2~q ),
	.datad(!\mii_rxdv_reg_2~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \packet_in_progress~0 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~1 (
	.dataa(!mii_clk_ena1),
	.datab(!packet_in_progress1),
	.datac(!\packet_in_progress~0_combout ),
	.datad(!\always2~0_combout ),
	.datae(!\always2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~1 .extended_lut = "off";
defparam \packet_in_progress~1 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \packet_in_progress~1 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_mii_tx_if (
	reset,
	mii_txd_int_0,
	mii_txd_int_1,
	mii_txd_int_2,
	mii_txd_int_3,
	mii_txerr_int1,
	mii_txdv_int1,
	tx_en_s_1,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	ethernet_mode,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mii_txd_int_0;
output 	mii_txd_int_1;
output 	mii_txd_int_2;
output 	mii_txd_int_3;
output 	mii_txerr_int1;
output 	mii_txdv_int1;
input 	tx_en_s_1;
input 	rd_14_4;
input 	rd_14_0;
input 	rd_14_5;
input 	rd_14_1;
input 	rd_14_6;
input 	rd_14_2;
input 	rd_14_7;
input 	rd_14_3;
input 	tx_err;
input 	ethernet_mode;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \mii_pos~0_combout ;
wire \mii_pos~q ;
wire \mii_txd_int~0_combout ;
wire \mii_txd_int~1_combout ;
wire \mii_txd_int~2_combout ;
wire \mii_txd_int~3_combout ;
wire \mii_txerr_int~0_combout ;
wire \mii_txdv_int~0_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_33 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(reset),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.ethernet_mode(ethernet_mode),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

dffeas \mii_txd_int[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_txd_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_txd_int_0),
	.prn(vcc));
defparam \mii_txd_int[0] .is_wysiwyg = "true";
defparam \mii_txd_int[0] .power_up = "low";

dffeas \mii_txd_int[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_txd_int~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_txd_int_1),
	.prn(vcc));
defparam \mii_txd_int[1] .is_wysiwyg = "true";
defparam \mii_txd_int[1] .power_up = "low";

dffeas \mii_txd_int[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_txd_int~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_txd_int_2),
	.prn(vcc));
defparam \mii_txd_int[2] .is_wysiwyg = "true";
defparam \mii_txd_int[2] .power_up = "low";

dffeas \mii_txd_int[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_txd_int~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_txd_int_3),
	.prn(vcc));
defparam \mii_txd_int[3] .is_wysiwyg = "true";
defparam \mii_txd_int[3] .power_up = "low";

dffeas mii_txerr_int(
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_txerr_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_txerr_int1),
	.prn(vcc));
defparam mii_txerr_int.is_wysiwyg = "true";
defparam mii_txerr_int.power_up = "low";

dffeas mii_txdv_int(
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_txdv_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mii_txdv_int1),
	.prn(vcc));
defparam mii_txdv_int.is_wysiwyg = "true";
defparam mii_txdv_int.power_up = "low";

cyclonev_lcell_comb \mii_pos~0 (
	.dataa(!tx_en_s_1),
	.datab(!\mii_pos~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_pos~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_pos~0 .extended_lut = "off";
defparam \mii_pos~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mii_pos~0 .shared_arith = "off";

dffeas mii_pos(
	.clk(mac_tx_clock_connection_clk),
	.d(\mii_pos~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mii_pos~q ),
	.prn(vcc));
defparam mii_pos.is_wysiwyg = "true";
defparam mii_pos.power_up = "low";

cyclonev_lcell_comb \mii_txd_int~0 (
	.dataa(!rd_14_4),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(!\mii_pos~q ),
	.datad(!rd_14_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_txd_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_txd_int~0 .extended_lut = "off";
defparam \mii_txd_int~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \mii_txd_int~0 .shared_arith = "off";

cyclonev_lcell_comb \mii_txd_int~1 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\mii_pos~q ),
	.datac(!rd_14_5),
	.datad(!rd_14_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_txd_int~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_txd_int~1 .extended_lut = "off";
defparam \mii_txd_int~1 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \mii_txd_int~1 .shared_arith = "off";

cyclonev_lcell_comb \mii_txd_int~2 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\mii_pos~q ),
	.datac(!rd_14_6),
	.datad(!rd_14_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_txd_int~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_txd_int~2 .extended_lut = "off";
defparam \mii_txd_int~2 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \mii_txd_int~2 .shared_arith = "off";

cyclonev_lcell_comb \mii_txd_int~3 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\mii_pos~q ),
	.datac(!rd_14_7),
	.datad(!rd_14_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_txd_int~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_txd_int~3 .extended_lut = "off";
defparam \mii_txd_int~3 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \mii_txd_int~3 .shared_arith = "off";

cyclonev_lcell_comb \mii_txerr_int~0 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!tx_err),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_txerr_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_txerr_int~0 .extended_lut = "off";
defparam \mii_txerr_int~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mii_txerr_int~0 .shared_arith = "off";

cyclonev_lcell_comb \mii_txdv_int~0 (
	.dataa(!tx_en_s_1),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mii_txdv_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mii_txdv_int~0 .extended_lut = "off";
defparam \mii_txdv_int~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mii_txdv_int~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_33 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	ethernet_mode,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	ethernet_mode;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_33 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(ethernet_mode),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_33 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_top_w_fifo (
	en,
	data_3,
	data_2,
	data_1,
	data_0,
	data_7,
	data_6,
	data_5,
	data_4,
	err,
	septy_flag,
	tx_ff_uflow,
	afull_flag,
	aempty_flag,
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	ff_rx_err_stat_5,
	ff_rx_err_stat_6,
	ff_rx_err_stat_7,
	ff_rx_err_stat_8,
	ff_rx_err_stat_9,
	ff_rx_err_stat_10,
	ff_rx_err_stat_11,
	ff_rx_err_stat_12,
	ff_rx_err_stat_13,
	ff_rx_err_stat_14,
	ff_rx_err_stat_15,
	ff_rx_err_stat_16,
	ff_rx_err_stat_17,
	ff_rx_err_stat_18,
	ff_rx_err_stat_19,
	ff_rx_err_stat_20,
	ff_rx_err_stat_4,
	ff_rx_err_stat_22,
	ff_rx_ucast,
	ff_rx_mcast,
	ff_rx_bcast,
	ff_rx_vlan,
	sav_flag,
	afull_flag1,
	aempty_flag1,
	altera_tse_reset_synchronizer_chain_out,
	txclk_ena,
	altera_tse_reset_synchronizer_chain_out1,
	altera_tse_reset_synchronizer_chain_out2,
	altera_tse_reset_synchronizer_chain_out3,
	tx_en_s_1,
	rxclk_ena,
	LessThan0,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	magic_detect,
	ethernet_mode,
	sleep_ena,
	dreg_1,
	m_rx_crs,
	dreg_11,
	din_s1,
	GND_port,
	clk_32_clk,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk,
	mac_misc_connection_ff_tx_crc_fwd)/* synthesis synthesis_greybox=1 */;
input 	en;
input 	data_3;
input 	data_2;
input 	data_1;
input 	data_0;
input 	data_7;
input 	data_6;
input 	data_5;
input 	data_4;
input 	err;
output 	septy_flag;
output 	tx_ff_uflow;
output 	afull_flag;
output 	aempty_flag;
output 	stateLOC_STATE_DATA;
output 	stateLOC_STATE_SHIFT;
output 	ff_rx_err_stat_5;
output 	ff_rx_err_stat_6;
output 	ff_rx_err_stat_7;
output 	ff_rx_err_stat_8;
output 	ff_rx_err_stat_9;
output 	ff_rx_err_stat_10;
output 	ff_rx_err_stat_11;
output 	ff_rx_err_stat_12;
output 	ff_rx_err_stat_13;
output 	ff_rx_err_stat_14;
output 	ff_rx_err_stat_15;
output 	ff_rx_err_stat_16;
output 	ff_rx_err_stat_17;
output 	ff_rx_err_stat_18;
output 	ff_rx_err_stat_19;
output 	ff_rx_err_stat_20;
output 	ff_rx_err_stat_4;
output 	ff_rx_err_stat_22;
output 	ff_rx_ucast;
output 	ff_rx_mcast;
output 	ff_rx_bcast;
output 	ff_rx_vlan;
output 	sav_flag;
output 	afull_flag1;
output 	aempty_flag1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	txclk_ena;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	altera_tse_reset_synchronizer_chain_out2;
input 	altera_tse_reset_synchronizer_chain_out3;
output 	tx_en_s_1;
input 	rxclk_ena;
input 	LessThan0;
output 	rd_14_4;
output 	rd_14_0;
output 	rd_14_5;
output 	rd_14_1;
output 	rd_14_6;
output 	rd_14_2;
output 	rd_14_7;
output 	rd_14_3;
output 	tx_err;
output 	magic_detect;
input 	ethernet_mode;
input 	sleep_ena;
input 	dreg_1;
input 	m_rx_crs;
input 	dreg_11;
output 	din_s1;
input 	GND_port;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;
input 	mac_misc_connection_ff_tx_crc_fwd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[9] ;
wire \U_TXFF|eop_sft[0]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[8] ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[4] ;
wire \U_TXFF|dout_reg_sft[28]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[0] ;
wire \U_TXFF|dout_reg_sft[24]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[5] ;
wire \U_TXFF|dout_reg_sft[29]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[1] ;
wire \U_TXFF|dout_reg_sft[25]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[6] ;
wire \U_TXFF|dout_reg_sft[30]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[2] ;
wire \U_TXFF|dout_reg_sft[26]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[7] ;
wire \U_TXFF|dout_reg_sft[31]~q ;
wire \U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[3] ;
wire \U_TXFF|dout_reg_sft[27]~q ;
wire \U_GETH|U_RX|rx_stat_wren~q ;
wire \U_GETH|U_RX|payload_length[0]~q ;
wire \U_GETH|U_RX|payload_length[1]~q ;
wire \U_GETH|U_RX|payload_length[2]~q ;
wire \U_GETH|U_RX|payload_length[3]~q ;
wire \U_GETH|U_RX|payload_length[4]~q ;
wire \U_GETH|U_RX|payload_length[5]~q ;
wire \U_GETH|U_RX|payload_length[6]~q ;
wire \U_GETH|U_RX|payload_length[7]~q ;
wire \U_GETH|U_RX|payload_length[8]~q ;
wire \U_GETH|U_RX|payload_length[9]~q ;
wire \U_GETH|U_RX|payload_length[10]~q ;
wire \U_GETH|U_RX|payload_length[11]~q ;
wire \U_GETH|U_RX|payload_length[12]~q ;
wire \U_GETH|U_RX|payload_length[13]~q ;
wire \U_GETH|U_RX|payload_length[14]~q ;
wire \U_GETH|U_RX|payload_length[15]~q ;
wire \U_TXFF|tx_empty~q ;
wire \U_TXFF|tx_data_int[7]~0_combout ;
wire \U_GETH|U_TX|U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \U_GETH|U_RX|rx_wren_int~q ;
wire \U_GETH|U_RX|rx_eop_int~q ;
wire \U_GETH|U_RX|rx_stat_data_s[5]~q ;
wire \U_GETH|U_RX|rx_stat_data_s[0]~q ;
wire \U_GETH|U_RX|rx_stat_data_s[1]~q ;
wire \U_GETH|U_RX|rx_stat_data_s[2]~q ;
wire \U_GETH|U_RX|rx_stat_data_s[3]~q ;
wire \U_GETH|U_RX|rx_sop_int~q ;
wire \U_GETH|U_RX|rx_ucast~q ;
wire \U_GETH|U_RX|rx_mcast~q ;
wire \U_GETH|U_RX|rx_bcast~q ;
wire \U_TXFF|tx_eop_int~0_combout ;
wire \U_TXFF|TX_STATUS|empty_flag~q ;
wire \U_GETH|U_TX|always9~1_combout ;
wire \U_GETH|U_TX|col_int~q ;
wire \U_GETH|U_TX|always9~3_combout ;
wire \U_GETH|U_TX|tx_rden_mii~q ;
wire \U_GETH|U_TX|tx_rden_int~0_combout ;
wire \U_GETH|U_TX|always9~4_combout ;
wire \U_TXFF|U_RETR|mac_ena~q ;
wire \U_TXFF|TX_DATA|sav_flag~q ;
wire \U_GETH|U_RX|rx_data_val~q ;
wire \U_GETH|U_RX|magic_pkt_ena~q ;
wire \U_GETH|U_TX|U_SYNC_6|std_sync_no_cut|dreg[1]~q ;
wire \U_TXFF|tx_stat[1]~q ;
wire \U_GETH|U_RX|rx_done_reg~q ;
wire \U_TXFF|sop_reg~q ;
wire \U_GETH|U_TX|tx_stat_rden~q ;
wire \U_GETH|U_RX|rx_data_int[3]~q ;
wire \U_GETH|U_RX|rx_data_int[2]~q ;
wire \U_GETH|U_RX|rx_data_int[1]~q ;
wire \U_GETH|U_RX|rx_data_int[0]~q ;
wire \U_GETH|U_RX|rx_data_int[7]~q ;
wire \U_GETH|U_RX|rx_data_int[6]~q ;
wire \U_GETH|U_RX|rx_data_int[5]~q ;
wire \U_GETH|U_RX|rx_data_int[4]~q ;
wire \U_TXFF|tx_stat[0]~q ;


IoTOctopus_QSYS_altera_tse_magic_detection U_MAGIC(
	.reset(altera_tse_reset_synchronizer_chain_out3),
	.clk_ena(rxclk_ena),
	.magic_detect1(magic_detect),
	.mac_data_val(\U_GETH|U_RX|rx_data_val~q ),
	.magic_pkt_ena(\U_GETH|U_RX|magic_pkt_ena~q ),
	.mac_data({\U_GETH|U_RX|rx_data_int[7]~q ,\U_GETH|U_RX|rx_data_int[6]~q ,\U_GETH|U_RX|rx_data_int[5]~q ,\U_GETH|U_RX|rx_data_int[4]~q ,\U_GETH|U_RX|rx_data_int[3]~q ,\U_GETH|U_RX|rx_data_int[2]~q ,\U_GETH|U_RX|rx_data_int[1]~q ,\U_GETH|U_RX|rx_data_int[0]~q }),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_top_1geth U_GETH(
	.q_b_9(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[9] ),
	.eop_sft_0(\U_TXFF|eop_sft[0]~q ),
	.q_b_8(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[8] ),
	.en(en),
	.data_3(data_3),
	.data_2(data_2),
	.data_1(data_1),
	.data_0(data_0),
	.data_7(data_7),
	.data_6(data_6),
	.data_5(data_5),
	.data_4(data_4),
	.q_b_4(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[4] ),
	.dout_reg_sft_28(\U_TXFF|dout_reg_sft[28]~q ),
	.q_b_0(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[0] ),
	.dout_reg_sft_24(\U_TXFF|dout_reg_sft[24]~q ),
	.q_b_5(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[5] ),
	.dout_reg_sft_29(\U_TXFF|dout_reg_sft[29]~q ),
	.q_b_1(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[1] ),
	.dout_reg_sft_25(\U_TXFF|dout_reg_sft[25]~q ),
	.q_b_6(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[6] ),
	.dout_reg_sft_30(\U_TXFF|dout_reg_sft[30]~q ),
	.q_b_2(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[2] ),
	.dout_reg_sft_26(\U_TXFF|dout_reg_sft[26]~q ),
	.q_b_7(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[7] ),
	.dout_reg_sft_31(\U_TXFF|dout_reg_sft[31]~q ),
	.q_b_3(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[3] ),
	.dout_reg_sft_27(\U_TXFF|dout_reg_sft[27]~q ),
	.err(err),
	.tx_ff_uflow(tx_ff_uflow),
	.afull_flag(afull_flag1),
	.txclk_ena(txclk_ena),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.rx_stat_wren(\U_GETH|U_RX|rx_stat_wren~q ),
	.payload_length_0(\U_GETH|U_RX|payload_length[0]~q ),
	.payload_length_1(\U_GETH|U_RX|payload_length[1]~q ),
	.payload_length_2(\U_GETH|U_RX|payload_length[2]~q ),
	.payload_length_3(\U_GETH|U_RX|payload_length[3]~q ),
	.payload_length_4(\U_GETH|U_RX|payload_length[4]~q ),
	.payload_length_5(\U_GETH|U_RX|payload_length[5]~q ),
	.payload_length_6(\U_GETH|U_RX|payload_length[6]~q ),
	.payload_length_7(\U_GETH|U_RX|payload_length[7]~q ),
	.payload_length_8(\U_GETH|U_RX|payload_length[8]~q ),
	.payload_length_9(\U_GETH|U_RX|payload_length[9]~q ),
	.payload_length_10(\U_GETH|U_RX|payload_length[10]~q ),
	.payload_length_11(\U_GETH|U_RX|payload_length[11]~q ),
	.payload_length_12(\U_GETH|U_RX|payload_length[12]~q ),
	.payload_length_13(\U_GETH|U_RX|payload_length[13]~q ),
	.payload_length_14(\U_GETH|U_RX|payload_length[14]~q ),
	.payload_length_15(\U_GETH|U_RX|payload_length[15]~q ),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out3),
	.tx_empty(\U_TXFF|tx_empty~q ),
	.tx_data_int_7(\U_TXFF|tx_data_int[7]~0_combout ),
	.dreg_1(\U_GETH|U_TX|U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.tx_en_s_1(tx_en_s_1),
	.rxclk_ena(rxclk_ena),
	.rx_wren_int(\U_GETH|U_RX|rx_wren_int~q ),
	.rx_eop_int(\U_GETH|U_RX|rx_eop_int~q ),
	.rx_stat_data_s_5(\U_GETH|U_RX|rx_stat_data_s[5]~q ),
	.rx_stat_data_s_0(\U_GETH|U_RX|rx_stat_data_s[0]~q ),
	.rx_stat_data_s_1(\U_GETH|U_RX|rx_stat_data_s[1]~q ),
	.rx_stat_data_s_2(\U_GETH|U_RX|rx_stat_data_s[2]~q ),
	.rx_stat_data_s_3(\U_GETH|U_RX|rx_stat_data_s[3]~q ),
	.rx_sop_int(\U_GETH|U_RX|rx_sop_int~q ),
	.rx_ucast(\U_GETH|U_RX|rx_ucast~q ),
	.rx_mcast(\U_GETH|U_RX|rx_mcast~q ),
	.rx_bcast(\U_GETH|U_RX|rx_bcast~q ),
	.rd_14_4(rd_14_4),
	.rd_14_0(rd_14_0),
	.rd_14_5(rd_14_5),
	.rd_14_1(rd_14_1),
	.rd_14_6(rd_14_6),
	.rd_14_2(rd_14_2),
	.rd_14_7(rd_14_7),
	.rd_14_3(rd_14_3),
	.tx_err(tx_err),
	.tx_eop_int(\U_TXFF|tx_eop_int~0_combout ),
	.empty_flag(\U_TXFF|TX_STATUS|empty_flag~q ),
	.always9(\U_GETH|U_TX|always9~1_combout ),
	.col_int(\U_GETH|U_TX|col_int~q ),
	.always91(\U_GETH|U_TX|always9~3_combout ),
	.tx_rden_mii(\U_GETH|U_TX|tx_rden_mii~q ),
	.tx_rden_int(\U_GETH|U_TX|tx_rden_int~0_combout ),
	.always92(\U_GETH|U_TX|always9~4_combout ),
	.mac_ena(\U_TXFF|U_RETR|mac_ena~q ),
	.sav_flag(\U_TXFF|TX_DATA|sav_flag~q ),
	.rx_data_val(\U_GETH|U_RX|rx_data_val~q ),
	.magic_pkt_ena(\U_GETH|U_RX|magic_pkt_ena~q ),
	.ethernet_mode(ethernet_mode),
	.dreg_11(\U_GETH|U_TX|U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.tx_stat_1(\U_TXFF|tx_stat[1]~q ),
	.rx_done_reg(\U_GETH|U_RX|rx_done_reg~q ),
	.sop_reg(\U_TXFF|sop_reg~q ),
	.tx_stat_rden(\U_GETH|U_TX|tx_stat_rden~q ),
	.sleep_ena(sleep_ena),
	.rx_data_int_3(\U_GETH|U_RX|rx_data_int[3]~q ),
	.rx_data_int_2(\U_GETH|U_RX|rx_data_int[2]~q ),
	.rx_data_int_1(\U_GETH|U_RX|rx_data_int[1]~q ),
	.rx_data_int_0(\U_GETH|U_RX|rx_data_int[0]~q ),
	.rx_data_int_7(\U_GETH|U_RX|rx_data_int[7]~q ),
	.rx_data_int_6(\U_GETH|U_RX|rx_data_int[6]~q ),
	.rx_data_int_5(\U_GETH|U_RX|rx_data_int[5]~q ),
	.rx_data_int_4(\U_GETH|U_RX|rx_data_int[4]~q ),
	.dreg_12(dreg_1),
	.m_rx_crs(m_rx_crs),
	.tx_stat_0(\U_TXFF|tx_stat[0]~q ),
	.GND_port(GND_port),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_rx_min_ff U_RXFF(
	.stateLOC_STATE_DATA(stateLOC_STATE_DATA),
	.stateLOC_STATE_SHIFT(stateLOC_STATE_SHIFT),
	.ff_rx_err_stat_5(ff_rx_err_stat_5),
	.ff_rx_err_stat_6(ff_rx_err_stat_6),
	.ff_rx_err_stat_7(ff_rx_err_stat_7),
	.ff_rx_err_stat_8(ff_rx_err_stat_8),
	.ff_rx_err_stat_9(ff_rx_err_stat_9),
	.ff_rx_err_stat_10(ff_rx_err_stat_10),
	.ff_rx_err_stat_11(ff_rx_err_stat_11),
	.ff_rx_err_stat_12(ff_rx_err_stat_12),
	.ff_rx_err_stat_13(ff_rx_err_stat_13),
	.ff_rx_err_stat_14(ff_rx_err_stat_14),
	.ff_rx_err_stat_15(ff_rx_err_stat_15),
	.ff_rx_err_stat_16(ff_rx_err_stat_16),
	.ff_rx_err_stat_17(ff_rx_err_stat_17),
	.ff_rx_err_stat_18(ff_rx_err_stat_18),
	.ff_rx_err_stat_19(ff_rx_err_stat_19),
	.ff_rx_err_stat_20(ff_rx_err_stat_20),
	.ff_rx_err_stat_4(ff_rx_err_stat_4),
	.ff_rx_err_stat_22(ff_rx_err_stat_22),
	.ff_rx_ucast(ff_rx_ucast),
	.ff_rx_mcast(ff_rx_mcast),
	.ff_rx_bcast(ff_rx_bcast),
	.ff_rx_vlan(ff_rx_vlan),
	.sav_flag(sav_flag),
	.afull_flag(afull_flag1),
	.aempty_flag(aempty_flag1),
	.rx_stat_wren(\U_GETH|U_RX|rx_stat_wren~q ),
	.payload_length_0(\U_GETH|U_RX|payload_length[0]~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out2),
	.payload_length_1(\U_GETH|U_RX|payload_length[1]~q ),
	.payload_length_2(\U_GETH|U_RX|payload_length[2]~q ),
	.payload_length_3(\U_GETH|U_RX|payload_length[3]~q ),
	.payload_length_4(\U_GETH|U_RX|payload_length[4]~q ),
	.payload_length_5(\U_GETH|U_RX|payload_length[5]~q ),
	.payload_length_6(\U_GETH|U_RX|payload_length[6]~q ),
	.payload_length_7(\U_GETH|U_RX|payload_length[7]~q ),
	.payload_length_8(\U_GETH|U_RX|payload_length[8]~q ),
	.payload_length_9(\U_GETH|U_RX|payload_length[9]~q ),
	.payload_length_10(\U_GETH|U_RX|payload_length[10]~q ),
	.payload_length_11(\U_GETH|U_RX|payload_length[11]~q ),
	.payload_length_12(\U_GETH|U_RX|payload_length[12]~q ),
	.payload_length_13(\U_GETH|U_RX|payload_length[13]~q ),
	.payload_length_14(\U_GETH|U_RX|payload_length[14]~q ),
	.payload_length_15(\U_GETH|U_RX|payload_length[15]~q ),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out3),
	.rx_wren_int(\U_GETH|U_RX|rx_wren_int~q ),
	.rx_eop_int(\U_GETH|U_RX|rx_eop_int~q ),
	.ff_rx_rdy(LessThan0),
	.rx_stat_data_s_5(\U_GETH|U_RX|rx_stat_data_s[5]~q ),
	.rx_stat_data_s_0(\U_GETH|U_RX|rx_stat_data_s[0]~q ),
	.rx_stat_data_s_1(\U_GETH|U_RX|rx_stat_data_s[1]~q ),
	.rx_stat_data_s_2(\U_GETH|U_RX|rx_stat_data_s[2]~q ),
	.rx_stat_data_s_3(\U_GETH|U_RX|rx_stat_data_s[3]~q ),
	.rx_sop_int(\U_GETH|U_RX|rx_sop_int~q ),
	.rx_ucast(\U_GETH|U_RX|rx_ucast~q ),
	.rx_mcast(\U_GETH|U_RX|rx_mcast~q ),
	.rx_bcast(\U_GETH|U_RX|rx_bcast~q ),
	.rx_done_reg(\U_GETH|U_RX|rx_done_reg~q ),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_tx_min_ff U_TXFF(
	.q_b_9(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[9] ),
	.eop_sft_0(\U_TXFF|eop_sft[0]~q ),
	.q_b_8(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[8] ),
	.q_b_4(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[4] ),
	.dout_reg_sft_28(\U_TXFF|dout_reg_sft[28]~q ),
	.q_b_0(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[0] ),
	.dout_reg_sft_24(\U_TXFF|dout_reg_sft[24]~q ),
	.q_b_5(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[5] ),
	.dout_reg_sft_29(\U_TXFF|dout_reg_sft[29]~q ),
	.q_b_1(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[1] ),
	.dout_reg_sft_25(\U_TXFF|dout_reg_sft[25]~q ),
	.q_b_6(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[6] ),
	.dout_reg_sft_30(\U_TXFF|dout_reg_sft[30]~q ),
	.q_b_2(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[2] ),
	.dout_reg_sft_26(\U_TXFF|dout_reg_sft[26]~q ),
	.q_b_7(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[7] ),
	.dout_reg_sft_31(\U_TXFF|dout_reg_sft[31]~q ),
	.q_b_3(\U_TXFF|U_RTSM|altsyncram_component|auto_generated|q_b[3] ),
	.dout_reg_sft_27(\U_TXFF|dout_reg_sft[27]~q ),
	.septy_flag(septy_flag),
	.afull_flag(afull_flag),
	.aempty_flag(aempty_flag),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.txclk_ena(txclk_ena),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.tx_empty1(\U_TXFF|tx_empty~q ),
	.tx_data_int_7(\U_TXFF|tx_data_int[7]~0_combout ),
	.dreg_1(\U_GETH|U_TX|U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.tx_eop_int(\U_TXFF|tx_eop_int~0_combout ),
	.empty_flag(\U_TXFF|TX_STATUS|empty_flag~q ),
	.always9(\U_GETH|U_TX|always9~1_combout ),
	.col_int(\U_GETH|U_TX|col_int~q ),
	.always91(\U_GETH|U_TX|always9~3_combout ),
	.tx_rden_mii(\U_GETH|U_TX|tx_rden_mii~q ),
	.tx_rden_int(\U_GETH|U_TX|tx_rden_int~0_combout ),
	.always92(\U_GETH|U_TX|always9~4_combout ),
	.mac_ena(\U_TXFF|U_RETR|mac_ena~q ),
	.sav_flag(\U_TXFF|TX_DATA|sav_flag~q ),
	.dreg_11(\U_GETH|U_TX|U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.tx_stat_1(\U_TXFF|tx_stat[1]~q ),
	.sop_reg1(\U_TXFF|sop_reg~q ),
	.tx_stat_rden(\U_GETH|U_TX|tx_stat_rden~q ),
	.dreg_12(dreg_11),
	.tx_stat_0(\U_TXFF|tx_stat[0]~q ),
	.din_s1(din_s1),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk),
	.mac_misc_connection_ff_tx_crc_fwd(mac_misc_connection_ff_tx_crc_fwd));

endmodule

module IoTOctopus_QSYS_altera_tse_magic_detection (
	reset,
	clk_ena,
	magic_detect1,
	mac_data_val,
	magic_pkt_ena,
	mac_data,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clk_ena;
output 	magic_detect1;
input 	mac_data_val;
input 	magic_pkt_ena;
input 	[7:0] mac_data;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \mac_data_val_reg~q ;
wire \mac_data_reg[3]~q ;
wire \mac_data_reg[2]~q ;
wire \mac_data_reg[1]~q ;
wire \mac_data_reg[0]~q ;
wire \mac_data_reg[7]~q ;
wire \mac_data_reg[6]~q ;
wire \mac_data_reg[5]~q ;
wire \mac_data_reg[4]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \addr_match1~q ;
wire \state~30_combout ;
wire \always3~0_combout ;
wire \always3~1_combout ;
wire \pbl_match~q ;
wire \Selector1~0_combout ;
wire \state~40_combout ;
wire \state.STM_TYP_IDLE~q ;
wire \Selector1~1_combout ;
wire \state~34_combout ;
wire \state.STM_TYP_WAIT_PBL~q ;
wire \pbl_cnt~3_combout ;
wire \pbl_cnt[0]~1_combout ;
wire \pbl_cnt[0]~q ;
wire \pbl_cnt~2_combout ;
wire \pbl_cnt[1]~q ;
wire \pbl_cnt~0_combout ;
wire \pbl_cnt[2]~q ;
wire \Equal8~0_combout ;
wire \pbl_cnt_dec~q ;
wire \state~41_combout ;
wire \state~42_combout ;
wire \state.STM_TYP_PBL~q ;
wire \state~36_combout ;
wire \state~37_combout ;
wire \state.STM_TYP_PAT0~q ;
wire \state~38_combout ;
wire \state.STM_TYP_PAT1~q ;
wire \state~39_combout ;
wire \state.STM_TYP_PAT2~q ;
wire \state~35_combout ;
wire \state.STM_TYP_PAT3~q ;
wire \state~33_combout ;
wire \state.STM_TYP_PAT4~q ;
wire \state~32_combout ;
wire \state.STM_TYP_PAT5~q ;
wire \pat_cnt~4_combout ;
wire \pat_cnt[0]~1_combout ;
wire \pat_cnt[0]~q ;
wire \pat_cnt~3_combout ;
wire \pat_cnt[1]~q ;
wire \pat_cnt~2_combout ;
wire \pat_cnt[2]~q ;
wire \pat_cnt~0_combout ;
wire \pat_cnt[3]~q ;
wire \Equal7~0_combout ;
wire \pat_cnt_dec~q ;
wire \state~31_combout ;
wire \state.STM_TYP_WAKE~q ;
wire \magic_detect~0_combout ;
wire \magic_detect~1_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_34 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(reset),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

dffeas magic_detect(
	.clk(mac_rx_clock_connection_clk),
	.d(\magic_detect~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(magic_detect1),
	.prn(vcc));
defparam magic_detect.is_wysiwyg = "true";
defparam magic_detect.power_up = "low";

dffeas mac_data_val_reg(
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data_val),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_val_reg~q ),
	.prn(vcc));
defparam mac_data_val_reg.is_wysiwyg = "true";
defparam mac_data_val_reg.power_up = "low";

dffeas \mac_data_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[3]~q ),
	.prn(vcc));
defparam \mac_data_reg[3] .is_wysiwyg = "true";
defparam \mac_data_reg[3] .power_up = "low";

dffeas \mac_data_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[2]~q ),
	.prn(vcc));
defparam \mac_data_reg[2] .is_wysiwyg = "true";
defparam \mac_data_reg[2] .power_up = "low";

dffeas \mac_data_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[1]~q ),
	.prn(vcc));
defparam \mac_data_reg[1] .is_wysiwyg = "true";
defparam \mac_data_reg[1] .power_up = "low";

dffeas \mac_data_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[0]~q ),
	.prn(vcc));
defparam \mac_data_reg[0] .is_wysiwyg = "true";
defparam \mac_data_reg[0] .power_up = "low";

dffeas \mac_data_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[7]~q ),
	.prn(vcc));
defparam \mac_data_reg[7] .is_wysiwyg = "true";
defparam \mac_data_reg[7] .power_up = "low";

dffeas \mac_data_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[6]~q ),
	.prn(vcc));
defparam \mac_data_reg[6] .is_wysiwyg = "true";
defparam \mac_data_reg[6] .power_up = "low";

dffeas \mac_data_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[5]~q ),
	.prn(vcc));
defparam \mac_data_reg[5] .is_wysiwyg = "true";
defparam \mac_data_reg[5] .power_up = "low";

dffeas \mac_data_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(mac_data[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\mac_data_reg[4]~q ),
	.prn(vcc));
defparam \mac_data_reg[4] .is_wysiwyg = "true";
defparam \mac_data_reg[4] .power_up = "low";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!\mac_data_reg[7]~q ),
	.datab(!\mac_data_reg[6]~q ),
	.datac(!\mac_data_reg[5]~q ),
	.datad(!\mac_data_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!\mac_data_reg[3]~q ),
	.datab(!\mac_data_reg[2]~q ),
	.datac(!\mac_data_reg[1]~q ),
	.datad(!\mac_data_reg[0]~q ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal1~1 .shared_arith = "off";

dffeas addr_match1(
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\addr_match1~q ),
	.prn(vcc));
defparam addr_match1.is_wysiwyg = "true";
defparam addr_match1.power_up = "low";

cyclonev_lcell_comb \state~30 (
	.dataa(!magic_pkt_ena),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~30 .extended_lut = "off";
defparam \state~30 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \state~30 .shared_arith = "off";

cyclonev_lcell_comb \always3~0 (
	.dataa(!\mac_data_val_reg~q ),
	.datab(!\mac_data_reg[7]~q ),
	.datac(!\mac_data_reg[6]~q ),
	.datad(!\mac_data_reg[5]~q ),
	.datae(!\mac_data_reg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \always3~0 .shared_arith = "off";

cyclonev_lcell_comb \always3~1 (
	.dataa(!\mac_data_reg[3]~q ),
	.datab(!\mac_data_reg[2]~q ),
	.datac(!\mac_data_reg[1]~q ),
	.datad(!\mac_data_reg[0]~q ),
	.datae(!\always3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~1 .extended_lut = "off";
defparam \always3~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \always3~1 .shared_arith = "off";

dffeas pbl_match(
	.clk(mac_rx_clock_connection_clk),
	.d(\always3~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\pbl_match~q ),
	.prn(vcc));
defparam pbl_match.is_wysiwyg = "true";
defparam pbl_match.power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\state.STM_TYP_PAT5~q ),
	.datab(!\state.STM_TYP_PAT4~q ),
	.datac(!\state.STM_TYP_PAT3~q ),
	.datad(!\state.STM_TYP_PAT0~q ),
	.datae(!\state.STM_TYP_PAT1~q ),
	.dataf(!\state.STM_TYP_PAT2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \state~40 (
	.dataa(!clk_ena),
	.datab(!\mac_data_val_reg~q ),
	.datac(!magic_pkt_ena),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYP_WAIT_PBL~q ),
	.dataf(!\state.STM_TYP_IDLE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~40 .extended_lut = "off";
defparam \state~40 .lut_mask = 64'hFF7FBF3FFFFFFFFF;
defparam \state~40 .shared_arith = "off";

dffeas \state.STM_TYP_IDLE (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~40_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_IDLE~q ),
	.prn(vcc));
defparam \state.STM_TYP_IDLE .is_wysiwyg = "true";
defparam \state.STM_TYP_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!\mac_data_val_reg~q ),
	.datab(!magic_pkt_ena),
	.datac(!\state.STM_TYP_WAIT_PBL~q ),
	.datad(!\state.STM_TYP_IDLE~q ),
	.datae(!\pbl_match~q ),
	.dataf(!\state.STM_TYP_PBL~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \state~34 (
	.dataa(!clk_ena),
	.datab(!\addr_match1~q ),
	.datac(!\state~30_combout ),
	.datad(!\state.STM_TYP_WAIT_PBL~q ),
	.datae(!\Selector1~0_combout ),
	.dataf(!\Selector1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~34 .extended_lut = "off";
defparam \state~34 .lut_mask = 64'hDFFF8FFFFFFFFFFF;
defparam \state~34 .shared_arith = "off";

dffeas \state.STM_TYP_WAIT_PBL (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~34_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_WAIT_PBL~q ),
	.prn(vcc));
defparam \state.STM_TYP_WAIT_PBL .is_wysiwyg = "true";
defparam \state.STM_TYP_WAIT_PBL .power_up = "low";

cyclonev_lcell_comb \pbl_cnt~3 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\state.STM_TYP_PBL~q ),
	.datac(!\pbl_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pbl_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pbl_cnt~3 .extended_lut = "off";
defparam \pbl_cnt~3 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \pbl_cnt~3 .shared_arith = "off";

cyclonev_lcell_comb \pbl_cnt[0]~1 (
	.dataa(!clk_ena),
	.datab(!\mac_data_val_reg~q ),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\state.STM_TYP_WAIT_PBL~q ),
	.datae(!\state.STM_TYP_IDLE~q ),
	.dataf(!\state.STM_TYP_PBL~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pbl_cnt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pbl_cnt[0]~1 .extended_lut = "off";
defparam \pbl_cnt[0]~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \pbl_cnt[0]~1 .shared_arith = "off";

dffeas \pbl_cnt[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pbl_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pbl_cnt[0]~1_combout ),
	.q(\pbl_cnt[0]~q ),
	.prn(vcc));
defparam \pbl_cnt[0] .is_wysiwyg = "true";
defparam \pbl_cnt[0] .power_up = "low";

cyclonev_lcell_comb \pbl_cnt~2 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\state.STM_TYP_PBL~q ),
	.datac(!\pbl_cnt[1]~q ),
	.datad(!\pbl_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pbl_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pbl_cnt~2 .extended_lut = "off";
defparam \pbl_cnt~2 .lut_mask = 64'hBFFBBFFBBFFBBFFB;
defparam \pbl_cnt~2 .shared_arith = "off";

dffeas \pbl_cnt[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pbl_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pbl_cnt[0]~1_combout ),
	.q(\pbl_cnt[1]~q ),
	.prn(vcc));
defparam \pbl_cnt[1] .is_wysiwyg = "true";
defparam \pbl_cnt[1] .power_up = "low";

cyclonev_lcell_comb \pbl_cnt~0 (
	.dataa(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datab(!\state.STM_TYP_PBL~q ),
	.datac(!\pbl_cnt[2]~q ),
	.datad(!\pbl_cnt[1]~q ),
	.datae(!\pbl_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pbl_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pbl_cnt~0 .extended_lut = "off";
defparam \pbl_cnt~0 .lut_mask = 64'hFBBFBFFBFBBFBFFB;
defparam \pbl_cnt~0 .shared_arith = "off";

dffeas \pbl_cnt[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pbl_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pbl_cnt[0]~1_combout ),
	.q(\pbl_cnt[2]~q ),
	.prn(vcc));
defparam \pbl_cnt[2] .is_wysiwyg = "true";
defparam \pbl_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Equal8~0 (
	.dataa(!\pbl_cnt[2]~q ),
	.datab(!\pbl_cnt[1]~q ),
	.datac(!\pbl_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal8~0 .extended_lut = "off";
defparam \Equal8~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Equal8~0 .shared_arith = "off";

dffeas pbl_cnt_dec(
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal8~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\pbl_cnt_dec~q ),
	.prn(vcc));
defparam pbl_cnt_dec.is_wysiwyg = "true";
defparam pbl_cnt_dec.power_up = "low";

cyclonev_lcell_comb \state~41 (
	.dataa(!clk_ena),
	.datab(!\mac_data_val_reg~q ),
	.datac(!\state.STM_TYP_WAIT_PBL~q ),
	.datad(!\pbl_match~q ),
	.datae(!\state.STM_TYP_PBL~q ),
	.dataf(!\pbl_cnt_dec~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~41 .extended_lut = "off";
defparam \state~41 .lut_mask = 64'hBFFFFFFF1FFFFFFF;
defparam \state~41 .shared_arith = "off";

cyclonev_lcell_comb \state~42 (
	.dataa(!\state~30_combout ),
	.datab(!\state~41_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~42 .extended_lut = "off";
defparam \state~42 .lut_mask = 64'h7777777777777777;
defparam \state~42 .shared_arith = "off";

dffeas \state.STM_TYP_PBL (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~42_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PBL~q ),
	.prn(vcc));
defparam \state.STM_TYP_PBL .is_wysiwyg = "true";
defparam \state.STM_TYP_PBL .power_up = "low";

cyclonev_lcell_comb \state~36 (
	.dataa(!\pat_cnt_dec~q ),
	.datab(!\addr_match1~q ),
	.datac(!\state.STM_TYP_PAT5~q ),
	.datad(!\pbl_match~q ),
	.datae(!\state.STM_TYP_PBL~q ),
	.dataf(!\pbl_cnt_dec~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~36 .extended_lut = "off";
defparam \state~36 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \state~36 .shared_arith = "off";

cyclonev_lcell_comb \state~37 (
	.dataa(!clk_ena),
	.datab(!\state~30_combout ),
	.datac(!\state.STM_TYP_PAT0~q ),
	.datad(!\state~36_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~37 .extended_lut = "off";
defparam \state~37 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \state~37 .shared_arith = "off";

dffeas \state.STM_TYP_PAT0 (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~37_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PAT0~q ),
	.prn(vcc));
defparam \state.STM_TYP_PAT0 .is_wysiwyg = "true";
defparam \state.STM_TYP_PAT0 .power_up = "low";

cyclonev_lcell_comb \state~38 (
	.dataa(!clk_ena),
	.datab(!magic_pkt_ena),
	.datac(!\addr_match1~q ),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYP_PAT0~q ),
	.dataf(!\state.STM_TYP_PAT1~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~38 .extended_lut = "off";
defparam \state~38 .lut_mask = 64'hBF1FFFFFFFFFFFFF;
defparam \state~38 .shared_arith = "off";

dffeas \state.STM_TYP_PAT1 (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~38_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PAT1~q ),
	.prn(vcc));
defparam \state.STM_TYP_PAT1 .is_wysiwyg = "true";
defparam \state.STM_TYP_PAT1 .power_up = "low";

cyclonev_lcell_comb \state~39 (
	.dataa(!clk_ena),
	.datab(!magic_pkt_ena),
	.datac(!\addr_match1~q ),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYP_PAT1~q ),
	.dataf(!\state.STM_TYP_PAT2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~39 .extended_lut = "off";
defparam \state~39 .lut_mask = 64'hBF1FFFFFFFFFFFFF;
defparam \state~39 .shared_arith = "off";

dffeas \state.STM_TYP_PAT2 (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~39_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PAT2~q ),
	.prn(vcc));
defparam \state.STM_TYP_PAT2 .is_wysiwyg = "true";
defparam \state.STM_TYP_PAT2 .power_up = "low";

cyclonev_lcell_comb \state~35 (
	.dataa(!clk_ena),
	.datab(!magic_pkt_ena),
	.datac(!\addr_match1~q ),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYP_PAT3~q ),
	.dataf(!\state.STM_TYP_PAT2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~35 .extended_lut = "off";
defparam \state~35 .lut_mask = 64'hBF1FFFFFFFFFFFFF;
defparam \state~35 .shared_arith = "off";

dffeas \state.STM_TYP_PAT3 (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~35_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PAT3~q ),
	.prn(vcc));
defparam \state.STM_TYP_PAT3 .is_wysiwyg = "true";
defparam \state.STM_TYP_PAT3 .power_up = "low";

cyclonev_lcell_comb \state~33 (
	.dataa(!clk_ena),
	.datab(!magic_pkt_ena),
	.datac(!\addr_match1~q ),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYP_PAT4~q ),
	.dataf(!\state.STM_TYP_PAT3~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~33 .extended_lut = "off";
defparam \state~33 .lut_mask = 64'hBF1FFFFFFFFFFFFF;
defparam \state~33 .shared_arith = "off";

dffeas \state.STM_TYP_PAT4 (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~33_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PAT4~q ),
	.prn(vcc));
defparam \state.STM_TYP_PAT4 .is_wysiwyg = "true";
defparam \state.STM_TYP_PAT4 .power_up = "low";

cyclonev_lcell_comb \state~32 (
	.dataa(!clk_ena),
	.datab(!magic_pkt_ena),
	.datac(!\addr_match1~q ),
	.datad(!\state.STM_TYP_PAT5~q ),
	.datae(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\state.STM_TYP_PAT4~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~32 .extended_lut = "off";
defparam \state~32 .lut_mask = 64'hBFFF1FFFFFFFFFFF;
defparam \state~32 .shared_arith = "off";

dffeas \state.STM_TYP_PAT5 (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~32_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_PAT5~q ),
	.prn(vcc));
defparam \state.STM_TYP_PAT5 .is_wysiwyg = "true";
defparam \state.STM_TYP_PAT5 .power_up = "low";

cyclonev_lcell_comb \pat_cnt~4 (
	.dataa(!\state.STM_TYP_PAT5~q ),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(!\pat_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pat_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pat_cnt~4 .extended_lut = "off";
defparam \pat_cnt~4 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \pat_cnt~4 .shared_arith = "off";

cyclonev_lcell_comb \pat_cnt[0]~1 (
	.dataa(!clk_ena),
	.datab(!\mac_data_val_reg~q ),
	.datac(!\state.STM_TYP_PAT5~q ),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\state.STM_TYP_WAIT_PBL~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pat_cnt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pat_cnt[0]~1 .extended_lut = "off";
defparam \pat_cnt[0]~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \pat_cnt[0]~1 .shared_arith = "off";

dffeas \pat_cnt[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pat_cnt~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pat_cnt[0]~1_combout ),
	.q(\pat_cnt[0]~q ),
	.prn(vcc));
defparam \pat_cnt[0] .is_wysiwyg = "true";
defparam \pat_cnt[0] .power_up = "low";

cyclonev_lcell_comb \pat_cnt~3 (
	.dataa(!\state.STM_TYP_PAT5~q ),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(!\pat_cnt[1]~q ),
	.datad(!\pat_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pat_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pat_cnt~3 .extended_lut = "off";
defparam \pat_cnt~3 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \pat_cnt~3 .shared_arith = "off";

dffeas \pat_cnt[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pat_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pat_cnt[0]~1_combout ),
	.q(\pat_cnt[1]~q ),
	.prn(vcc));
defparam \pat_cnt[1] .is_wysiwyg = "true";
defparam \pat_cnt[1] .power_up = "low";

cyclonev_lcell_comb \pat_cnt~2 (
	.dataa(!\state.STM_TYP_PAT5~q ),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(!\pat_cnt[2]~q ),
	.datad(!\pat_cnt[1]~q ),
	.datae(!\pat_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pat_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pat_cnt~2 .extended_lut = "off";
defparam \pat_cnt~2 .lut_mask = 64'hFDDFDFFDFDDFDFFD;
defparam \pat_cnt~2 .shared_arith = "off";

dffeas \pat_cnt[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pat_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pat_cnt[0]~1_combout ),
	.q(\pat_cnt[2]~q ),
	.prn(vcc));
defparam \pat_cnt[2] .is_wysiwyg = "true";
defparam \pat_cnt[2] .power_up = "low";

cyclonev_lcell_comb \pat_cnt~0 (
	.dataa(!\state.STM_TYP_PAT5~q ),
	.datab(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datac(!\pat_cnt[3]~q ),
	.datad(!\pat_cnt[2]~q ),
	.datae(!\pat_cnt[1]~q ),
	.dataf(!\pat_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pat_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pat_cnt~0 .extended_lut = "off";
defparam \pat_cnt~0 .lut_mask = 64'hDFFDFDDFFDDFDFFD;
defparam \pat_cnt~0 .shared_arith = "off";

dffeas \pat_cnt[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\pat_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pat_cnt[0]~1_combout ),
	.q(\pat_cnt[3]~q ),
	.prn(vcc));
defparam \pat_cnt[3] .is_wysiwyg = "true";
defparam \pat_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Equal7~0 (
	.dataa(!\pat_cnt[3]~q ),
	.datab(!\pat_cnt[2]~q ),
	.datac(!\pat_cnt[1]~q ),
	.datad(!\pat_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal7~0 .extended_lut = "off";
defparam \Equal7~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal7~0 .shared_arith = "off";

dffeas pat_cnt_dec(
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal7~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\pat_cnt_dec~q ),
	.prn(vcc));
defparam pat_cnt_dec.is_wysiwyg = "true";
defparam pat_cnt_dec.power_up = "low";

cyclonev_lcell_comb \state~31 (
	.dataa(!clk_ena),
	.datab(!\state.STM_TYP_WAKE~q ),
	.datac(!\pat_cnt_dec~q ),
	.datad(!\addr_match1~q ),
	.datae(!\state.STM_TYP_PAT5~q ),
	.dataf(!\state~30_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~31 .extended_lut = "off";
defparam \state~31 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \state~31 .shared_arith = "off";

dffeas \state.STM_TYP_WAKE (
	.clk(mac_rx_clock_connection_clk),
	.d(\state~31_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_WAKE~q ),
	.prn(vcc));
defparam \state.STM_TYP_WAKE .is_wysiwyg = "true";
defparam \state.STM_TYP_WAKE .power_up = "low";

cyclonev_lcell_comb \magic_detect~0 (
	.dataa(!magic_pkt_ena),
	.datab(!\state.STM_TYP_WAKE~q ),
	.datac(!\pat_cnt_dec~q ),
	.datad(!\addr_match1~q ),
	.datae(!\state.STM_TYP_PAT5~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\magic_detect~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \magic_detect~0 .extended_lut = "off";
defparam \magic_detect~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \magic_detect~0 .shared_arith = "off";

cyclonev_lcell_comb \magic_detect~1 (
	.dataa(!magic_detect1),
	.datab(!mac_data_val),
	.datac(!\mac_data_val_reg~q ),
	.datad(!\magic_detect~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\magic_detect~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \magic_detect~1 .extended_lut = "off";
defparam \magic_detect~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \magic_detect~1 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_34 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_34 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_34 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_rx_min_ff (
	stateLOC_STATE_DATA,
	stateLOC_STATE_SHIFT,
	ff_rx_err_stat_5,
	ff_rx_err_stat_6,
	ff_rx_err_stat_7,
	ff_rx_err_stat_8,
	ff_rx_err_stat_9,
	ff_rx_err_stat_10,
	ff_rx_err_stat_11,
	ff_rx_err_stat_12,
	ff_rx_err_stat_13,
	ff_rx_err_stat_14,
	ff_rx_err_stat_15,
	ff_rx_err_stat_16,
	ff_rx_err_stat_17,
	ff_rx_err_stat_18,
	ff_rx_err_stat_19,
	ff_rx_err_stat_20,
	ff_rx_err_stat_4,
	ff_rx_err_stat_22,
	ff_rx_ucast,
	ff_rx_mcast,
	ff_rx_bcast,
	ff_rx_vlan,
	sav_flag,
	afull_flag,
	aempty_flag,
	rx_stat_wren,
	payload_length_0,
	altera_tse_reset_synchronizer_chain_out,
	payload_length_1,
	payload_length_2,
	payload_length_3,
	payload_length_4,
	payload_length_5,
	payload_length_6,
	payload_length_7,
	payload_length_8,
	payload_length_9,
	payload_length_10,
	payload_length_11,
	payload_length_12,
	payload_length_13,
	payload_length_14,
	payload_length_15,
	altera_tse_reset_synchronizer_chain_out1,
	rx_wren_int,
	rx_eop_int,
	ff_rx_rdy,
	rx_stat_data_s_5,
	rx_stat_data_s_0,
	rx_stat_data_s_1,
	rx_stat_data_s_2,
	rx_stat_data_s_3,
	rx_sop_int,
	rx_ucast,
	rx_mcast,
	rx_bcast,
	rx_done_reg,
	GND_port,
	clk_32_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	stateLOC_STATE_DATA;
output 	stateLOC_STATE_SHIFT;
output 	ff_rx_err_stat_5;
output 	ff_rx_err_stat_6;
output 	ff_rx_err_stat_7;
output 	ff_rx_err_stat_8;
output 	ff_rx_err_stat_9;
output 	ff_rx_err_stat_10;
output 	ff_rx_err_stat_11;
output 	ff_rx_err_stat_12;
output 	ff_rx_err_stat_13;
output 	ff_rx_err_stat_14;
output 	ff_rx_err_stat_15;
output 	ff_rx_err_stat_16;
output 	ff_rx_err_stat_17;
output 	ff_rx_err_stat_18;
output 	ff_rx_err_stat_19;
output 	ff_rx_err_stat_20;
output 	ff_rx_err_stat_4;
output 	ff_rx_err_stat_22;
output 	ff_rx_ucast;
output 	ff_rx_mcast;
output 	ff_rx_bcast;
output 	ff_rx_vlan;
output 	sav_flag;
output 	afull_flag;
output 	aempty_flag;
input 	rx_stat_wren;
input 	payload_length_0;
input 	altera_tse_reset_synchronizer_chain_out;
input 	payload_length_1;
input 	payload_length_2;
input 	payload_length_3;
input 	payload_length_4;
input 	payload_length_5;
input 	payload_length_6;
input 	payload_length_7;
input 	payload_length_8;
input 	payload_length_9;
input 	payload_length_10;
input 	payload_length_11;
input 	payload_length_12;
input 	payload_length_13;
input 	payload_length_14;
input 	payload_length_15;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	rx_wren_int;
input 	rx_eop_int;
input 	ff_rx_rdy;
input 	rx_stat_data_s_5;
input 	rx_stat_data_s_0;
input 	rx_stat_data_s_1;
input 	rx_stat_data_s_2;
input 	rx_stat_data_s_3;
input 	rx_sop_int;
input 	rx_ucast;
input 	rx_mcast;
input 	rx_bcast;
input 	rx_done_reg;
input 	GND_port;
input 	clk_32_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[5] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[6] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[7] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[8] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[9] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[10] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[11] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[12] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[13] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[14] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[15] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[16] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[17] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[18] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[19] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[20] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[4] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[22] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[36] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ;
wire \RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[37] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[21] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[2] ;
wire \RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[3] ;
wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \RX_STATUS|empty_flag~q ;
wire \rx_wren32~q ;
wire \rx_eop32~q ;
wire \U_SYNC_5|std_sync_no_cut|dreg[1]~q ;
wire \byte_empty[1]~q ;
wire \frm_type32[0]~q ;
wire \rx_sop32~q ;
wire \frm_type32[2]~q ;
wire \frm_type32[1]~q ;
wire \U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \byte_empty[0]~q ;
wire \always6~0_combout ;
wire \always4~0_combout ;
wire \data_rdreq~combout ;
wire \U_SYNC_4|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_6|std_sync_no_cut|dreg[1]~q ;
wire \byte_empty~0_combout ;
wire \byte_empty[0]~1_combout ;
wire \frm_type32~0_combout ;
wire \frm_type32[1]~1_combout ;
wire \rx_sop32~0_combout ;
wire \frm_type32~2_combout ;
wire \frm_type32~3_combout ;
wire \byte_empty~2_combout ;
wire \rx_rdy_reg~q ;
wire \Selector1~0_combout ;
wire \always10~0_combout ;
wire \Selector1~3_combout ;
wire \sw_reset_ff_flush~0_combout ;
wire \sw_reset_ff_flush_counter[0]~4_combout ;
wire \sw_reset_ff_flush_counter[0]~q ;
wire \sw_reset_ff_flush_counter[1]~3_combout ;
wire \sw_reset_ff_flush_counter[1]~q ;
wire \sw_reset_ff_flush~3_combout ;
wire \sw_reset_ff_flush_counter[2]~2_combout ;
wire \sw_reset_ff_flush_counter[2]~q ;
wire \sw_reset_ff_flush_counter[3]~1_combout ;
wire \sw_reset_ff_flush_counter[3]~q ;
wire \sw_reset_ff_flush~1_combout ;
wire \sw_reset_ff_flush_counter[4]~0_combout ;
wire \sw_reset_ff_flush_counter[4]~q ;
wire \sw_reset_ff_flush~2_combout ;
wire \sw_reset_ff_flush~q ;
wire \Selector2~0_combout ;
wire \state.LOC_STATE_WAIT~q ;
wire \always10~1_combout ;
wire \Selector0~0_combout ;
wire \Selector5~0_combout ;
wire \Selector9~0_combout ;
wire \state.LOC_STATE_FF_DATA_FLUSH_WAIT~q ;
wire \Selector5~1_combout ;
wire \Selector5~2_combout ;
wire \state.LOC_STATE_FF_DATA_FLUSH~q ;
wire \Selector6~0_combout ;
wire \state.LOC_STATE_FF_FLUSH_WAIT~q ;
wire \Selector4~0_combout ;
wire \Selector4~2_combout ;
wire \state.LOC_STATE_END_FRM~q ;
wire \Selector8~0_combout ;
wire \state.LOC_STATE_RST_DONE~q ;
wire \Selector0~1_combout ;
wire \Selector0~2_combout ;
wire \state.LOC_STATE_IDLE~q ;
wire \rx_err_sig~0_combout ;
wire \Selector1~1_combout ;
wire \Selector1~2_combout ;
wire \Selector7~0_combout ;
wire \state.LOC_STATE_SHIFT_WAIT~q ;
wire \Selector3~0_combout ;
wire \rx_frm_type_reg~0_combout ;
wire \Selector4~1_combout ;
wire \rx_frm_type_reg[1]~1_combout ;
wire \rx_frm_type_reg[0]~q ;
wire \rx_frm_type_reg~2_combout ;
wire \rx_frm_type_reg[2]~q ;
wire \rx_frm_type_reg~3_combout ;
wire \rx_frm_type_reg[1]~q ;
wire \rx_frm_type_reg~4_combout ;
wire \rx_frm_type_reg[3]~q ;


IoTOctopus_QSYS_altera_tse_a_fifo_34 RX_STATUS(
	.q_b_5(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[5] ),
	.q_b_6(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[6] ),
	.q_b_7(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[7] ),
	.q_b_8(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[8] ),
	.q_b_9(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[9] ),
	.q_b_10(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[10] ),
	.q_b_11(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[11] ),
	.q_b_12(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[12] ),
	.q_b_13(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[13] ),
	.q_b_14(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[14] ),
	.q_b_15(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[15] ),
	.q_b_16(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[16] ),
	.q_b_17(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[17] ),
	.q_b_18(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[18] ),
	.q_b_19(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[19] ),
	.q_b_20(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[20] ),
	.q_b_4(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[4] ),
	.q_b_22(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[22] ),
	.q_b_21(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[21] ),
	.q_b_0(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.q_b_1(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.q_b_2(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.q_b_3(\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.empty_flag1(\RX_STATUS|empty_flag~q ),
	.Selector4(\Selector4~0_combout ),
	.rx_stat_wren(rx_stat_wren),
	.payload_length_0(payload_length_0),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.Selector41(\Selector4~1_combout ),
	.payload_length_1(payload_length_1),
	.payload_length_2(payload_length_2),
	.payload_length_3(payload_length_3),
	.payload_length_4(payload_length_4),
	.payload_length_5(payload_length_5),
	.payload_length_6(payload_length_6),
	.payload_length_7(payload_length_7),
	.payload_length_8(payload_length_8),
	.payload_length_9(payload_length_9),
	.payload_length_10(payload_length_10),
	.payload_length_11(payload_length_11),
	.payload_length_12(payload_length_12),
	.payload_length_13(payload_length_13),
	.payload_length_14(payload_length_14),
	.payload_length_15(payload_length_15),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.Selector42(\Selector4~2_combout ),
	.rx_stat_data_s_5(rx_stat_data_s_5),
	.rx_stat_data_s_0(rx_stat_data_s_0),
	.rx_stat_data_s_1(rx_stat_data_s_1),
	.rx_stat_data_s_2(rx_stat_data_s_2),
	.rx_stat_data_s_3(rx_stat_data_s_3),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_a_fifo_opt_1246 RX_DATA(
	.q_b_32(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.q_b_39(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.q_b_34(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.q_b_33(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.q_b_36(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[36] ),
	.q_b_35(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.q_b_37(\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[37] ),
	.sav_flag1(sav_flag),
	.afull_flag1(afull_flag),
	.aempty_flag1(aempty_flag),
	.rx_wren32(\rx_wren32~q ),
	.rx_eop32(\rx_eop32~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.byte_empty_1(\byte_empty[1]~q ),
	.frm_type32_0(\frm_type32[0]~q ),
	.rx_sop32(\rx_sop32~q ),
	.frm_type32_2(\frm_type32[2]~q ),
	.frm_type32_1(\frm_type32[1]~q ),
	.dreg_1(\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.data_rdreq(\data_rdreq~combout ),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_38 U_SYNC_6(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.rx_done_reg(rx_done_reg),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_37 U_SYNC_5(
	.dreg_1(\U_SYNC_5|std_sync_no_cut|dreg[1]~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_36 U_SYNC_4(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_2 U_SYNC_2(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_35 U_SYNC_1(
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

dffeas rx_wren32(
	.clk(mac_rx_clock_connection_clk),
	.d(\always6~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rx_wren32~q ),
	.prn(vcc));
defparam rx_wren32.is_wysiwyg = "true";
defparam rx_wren32.power_up = "low";

dffeas rx_eop32(
	.clk(mac_rx_clock_connection_clk),
	.d(\always4~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rx_eop32~q ),
	.prn(vcc));
defparam rx_eop32.is_wysiwyg = "true";
defparam rx_eop32.power_up = "low";

dffeas \byte_empty[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\byte_empty~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\byte_empty[0]~1_combout ),
	.q(\byte_empty[1]~q ),
	.prn(vcc));
defparam \byte_empty[1] .is_wysiwyg = "true";
defparam \byte_empty[1] .power_up = "low";

dffeas \frm_type32[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_type32~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\frm_type32[1]~1_combout ),
	.q(\frm_type32[0]~q ),
	.prn(vcc));
defparam \frm_type32[0] .is_wysiwyg = "true";
defparam \frm_type32[0] .power_up = "low";

dffeas rx_sop32(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_sop32~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rx_sop32~q ),
	.prn(vcc));
defparam rx_sop32.is_wysiwyg = "true";
defparam rx_sop32.power_up = "low";

dffeas \frm_type32[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_type32~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\frm_type32[1]~1_combout ),
	.q(\frm_type32[2]~q ),
	.prn(vcc));
defparam \frm_type32[2] .is_wysiwyg = "true";
defparam \frm_type32[2] .power_up = "low";

dffeas \frm_type32[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_type32~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\frm_type32[1]~1_combout ),
	.q(\frm_type32[1]~q ),
	.prn(vcc));
defparam \frm_type32[1] .is_wysiwyg = "true";
defparam \frm_type32[1] .power_up = "low";

dffeas \byte_empty[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\byte_empty~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\byte_empty[0]~1_combout ),
	.q(\byte_empty[0]~q ),
	.prn(vcc));
defparam \byte_empty[0] .is_wysiwyg = "true";
defparam \byte_empty[0] .power_up = "low";

cyclonev_lcell_comb \always6~0 (
	.dataa(!\byte_empty[1]~q ),
	.datab(!rx_wren_int),
	.datac(!rx_eop_int),
	.datad(!\byte_empty[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \always6~0 .shared_arith = "off";

cyclonev_lcell_comb \always4~0 (
	.dataa(!rx_wren_int),
	.datab(!rx_eop_int),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'h7777777777777777;
defparam \always4~0 .shared_arith = "off";

cyclonev_lcell_comb data_rdreq(
	.dataa(!\Selector1~0_combout ),
	.datab(!\always10~0_combout ),
	.datac(!\state.LOC_STATE_WAIT~q ),
	.datad(!\sw_reset_ff_flush~q ),
	.datae(!\Selector1~1_combout ),
	.dataf(!\Selector5~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_rdreq~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam data_rdreq.extended_lut = "off";
defparam data_rdreq.lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam data_rdreq.shared_arith = "off";

cyclonev_lcell_comb \byte_empty~0 (
	.dataa(!\rx_eop32~q ),
	.datab(!\byte_empty[1]~q ),
	.datac(!rx_wren_int),
	.datad(!\byte_empty[0]~q ),
	.datae(!rx_sop_int),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_empty~0 .extended_lut = "off";
defparam \byte_empty~0 .lut_mask = 64'hBFEFFFFFBFEFFFFF;
defparam \byte_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \byte_empty[0]~1 (
	.dataa(!\rx_eop32~q ),
	.datab(!rx_wren_int),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_empty[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_empty[0]~1 .extended_lut = "off";
defparam \byte_empty[0]~1 .lut_mask = 64'h7777777777777777;
defparam \byte_empty[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \frm_type32~0 (
	.dataa(!rx_wren_int),
	.datab(!rx_sop_int),
	.datac(!rx_ucast),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_type32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_type32~0 .extended_lut = "off";
defparam \frm_type32~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \frm_type32~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_type32[1]~1 (
	.dataa(!\byte_empty[1]~q ),
	.datab(!rx_wren_int),
	.datac(!\byte_empty[0]~q ),
	.datad(!rx_sop_int),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_type32[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_type32[1]~1 .extended_lut = "off";
defparam \frm_type32[1]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \frm_type32[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rx_sop32~0 (
	.dataa(!\byte_empty[1]~q ),
	.datab(!\rx_sop32~q ),
	.datac(!rx_wren_int),
	.datad(!\byte_empty[0]~q ),
	.datae(!rx_sop_int),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_sop32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_sop32~0 .extended_lut = "off";
defparam \rx_sop32~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \rx_sop32~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_type32~2 (
	.dataa(!rx_wren_int),
	.datab(!rx_sop_int),
	.datac(!rx_mcast),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_type32~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_type32~2 .extended_lut = "off";
defparam \frm_type32~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \frm_type32~2 .shared_arith = "off";

cyclonev_lcell_comb \frm_type32~3 (
	.dataa(!rx_wren_int),
	.datab(!rx_sop_int),
	.datac(!rx_bcast),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_type32~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_type32~3 .extended_lut = "off";
defparam \frm_type32~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \frm_type32~3 .shared_arith = "off";

cyclonev_lcell_comb \byte_empty~2 (
	.dataa(!\rx_eop32~q ),
	.datab(!rx_wren_int),
	.datac(!\byte_empty[0]~q ),
	.datad(!rx_sop_int),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_empty~2 .extended_lut = "off";
defparam \byte_empty~2 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \byte_empty~2 .shared_arith = "off";

dffeas \state.LOC_STATE_DATA (
	.clk(clk_32_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateLOC_STATE_DATA),
	.prn(vcc));
defparam \state.LOC_STATE_DATA .is_wysiwyg = "true";
defparam \state.LOC_STATE_DATA .power_up = "low";

dffeas \state.LOC_STATE_SHIFT (
	.clk(clk_32_clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateLOC_STATE_SHIFT),
	.prn(vcc));
defparam \state.LOC_STATE_SHIFT .is_wysiwyg = "true";
defparam \state.LOC_STATE_SHIFT .power_up = "low";

cyclonev_lcell_comb \ff_rx_err_stat[5]~0 (
	.dataa(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[5] ),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datac(!stateLOC_STATE_DATA),
	.datad(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datae(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.dataf(!\Selector4~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[5]~0 .extended_lut = "off";
defparam \ff_rx_err_stat[5]~0 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \ff_rx_err_stat[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[6]~1 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[6] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[6]~1 .extended_lut = "off";
defparam \ff_rx_err_stat[6]~1 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[7]~2 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[7] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[7]~2 .extended_lut = "off";
defparam \ff_rx_err_stat[7]~2 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[7]~2 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[8]~3 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[8] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[8]~3 .extended_lut = "off";
defparam \ff_rx_err_stat[8]~3 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[8]~3 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[9]~4 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[9] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[9]~4 .extended_lut = "off";
defparam \ff_rx_err_stat[9]~4 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[9]~4 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[10]~5 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[10] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[10]~5 .extended_lut = "off";
defparam \ff_rx_err_stat[10]~5 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[10]~5 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[11]~6 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[11] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[11]~6 .extended_lut = "off";
defparam \ff_rx_err_stat[11]~6 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[11]~6 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[12]~7 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[12] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[12]~7 .extended_lut = "off";
defparam \ff_rx_err_stat[12]~7 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[12]~7 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[13]~8 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[13] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[13]~8 .extended_lut = "off";
defparam \ff_rx_err_stat[13]~8 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[13]~8 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[14]~9 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[14] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[14]~9 .extended_lut = "off";
defparam \ff_rx_err_stat[14]~9 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[14]~9 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[15]~10 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[15] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[15]~10 .extended_lut = "off";
defparam \ff_rx_err_stat[15]~10 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[15]~10 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[16]~11 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[16] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[16]~11 .extended_lut = "off";
defparam \ff_rx_err_stat[16]~11 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[16]~11 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[17]~12 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[17] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[17]~12 .extended_lut = "off";
defparam \ff_rx_err_stat[17]~12 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[17]~12 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[18]~13 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[18] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[18]~13 .extended_lut = "off";
defparam \ff_rx_err_stat[18]~13 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[18]~13 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[19]~14 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[19] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[19]~14 .extended_lut = "off";
defparam \ff_rx_err_stat[19]~14 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[19]~14 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[20]~15 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[20] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[20]~15 .extended_lut = "off";
defparam \ff_rx_err_stat[20]~15 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[20]~15 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[4]~16 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[4] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[4]~16 .extended_lut = "off";
defparam \ff_rx_err_stat[4]~16 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[4]~16 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_err_stat[22]~17 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[22] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_err_stat_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_err_stat[22]~17 .extended_lut = "off";
defparam \ff_rx_err_stat[22]~17 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \ff_rx_err_stat[22]~17 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_ucast~0 (
	.dataa(!stateLOC_STATE_DATA),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.datac(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datad(!\rx_frm_type_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_ucast),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_ucast~0 .extended_lut = "off";
defparam \ff_rx_ucast~0 .lut_mask = 64'h7BFF7BFF7BFF7BFF;
defparam \ff_rx_ucast~0 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_mcast~0 (
	.dataa(!stateLOC_STATE_DATA),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[36] ),
	.datad(!\rx_frm_type_reg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_mcast),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_mcast~0 .extended_lut = "off";
defparam \ff_rx_mcast~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ff_rx_mcast~0 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_bcast~0 (
	.dataa(!stateLOC_STATE_DATA),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.datad(!\rx_frm_type_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_bcast),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_bcast~0 .extended_lut = "off";
defparam \ff_rx_bcast~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ff_rx_bcast~0 .shared_arith = "off";

cyclonev_lcell_comb \ff_rx_vlan~0 (
	.dataa(!stateLOC_STATE_DATA),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[37] ),
	.datad(!\rx_frm_type_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(ff_rx_vlan),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rx_vlan~0 .extended_lut = "off";
defparam \ff_rx_vlan~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \ff_rx_vlan~0 .shared_arith = "off";

dffeas rx_rdy_reg(
	.clk(clk_32_clk),
	.d(ff_rx_rdy),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rx_rdy_reg~q ),
	.prn(vcc));
defparam rx_rdy_reg.is_wysiwyg = "true";
defparam rx_rdy_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datac(!stateLOC_STATE_DATA),
	.datad(!aempty_flag),
	.datae(!\rx_rdy_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!sav_flag),
	.datac(!\rx_rdy_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!aempty_flag),
	.datac(!\rx_rdy_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \sw_reset_ff_flush~0 (
	.dataa(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush~0 .extended_lut = "off";
defparam \sw_reset_ff_flush~0 .lut_mask = 64'h7777777777777777;
defparam \sw_reset_ff_flush~0 .shared_arith = "off";

cyclonev_lcell_comb \sw_reset_ff_flush_counter[0]~4 (
	.dataa(!\sw_reset_ff_flush_counter[4]~q ),
	.datab(!\sw_reset_ff_flush~0_combout ),
	.datac(!\sw_reset_ff_flush_counter[0]~q ),
	.datad(!\sw_reset_ff_flush~1_combout ),
	.datae(!ff_rx_rdy),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush_counter[0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush_counter[0]~4 .extended_lut = "off";
defparam \sw_reset_ff_flush_counter[0]~4 .lut_mask = 64'hF7FF37FFF7FF37FF;
defparam \sw_reset_ff_flush_counter[0]~4 .shared_arith = "off";

dffeas \sw_reset_ff_flush_counter[0] (
	.clk(clk_32_clk),
	.d(\sw_reset_ff_flush_counter[0]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sw_reset_ff_flush_counter[0]~q ),
	.prn(vcc));
defparam \sw_reset_ff_flush_counter[0] .is_wysiwyg = "true";
defparam \sw_reset_ff_flush_counter[0] .power_up = "low";

cyclonev_lcell_comb \sw_reset_ff_flush_counter[1]~3 (
	.dataa(!\sw_reset_ff_flush_counter[4]~q ),
	.datab(!\sw_reset_ff_flush~0_combout ),
	.datac(!\sw_reset_ff_flush_counter[1]~q ),
	.datad(!\sw_reset_ff_flush_counter[0]~q ),
	.datae(!\sw_reset_ff_flush~1_combout ),
	.dataf(!ff_rx_rdy),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush_counter[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush_counter[1]~3 .extended_lut = "off";
defparam \sw_reset_ff_flush_counter[1]~3 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \sw_reset_ff_flush_counter[1]~3 .shared_arith = "off";

dffeas \sw_reset_ff_flush_counter[1] (
	.clk(clk_32_clk),
	.d(\sw_reset_ff_flush_counter[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sw_reset_ff_flush_counter[1]~q ),
	.prn(vcc));
defparam \sw_reset_ff_flush_counter[1] .is_wysiwyg = "true";
defparam \sw_reset_ff_flush_counter[1] .power_up = "low";

cyclonev_lcell_comb \sw_reset_ff_flush~3 (
	.dataa(!\sw_reset_ff_flush_counter[1]~q ),
	.datab(!\sw_reset_ff_flush_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush~3 .extended_lut = "off";
defparam \sw_reset_ff_flush~3 .lut_mask = 64'h7777777777777777;
defparam \sw_reset_ff_flush~3 .shared_arith = "off";

cyclonev_lcell_comb \sw_reset_ff_flush_counter[2]~2 (
	.dataa(!\sw_reset_ff_flush_counter[4]~q ),
	.datab(!\sw_reset_ff_flush~0_combout ),
	.datac(!\sw_reset_ff_flush_counter[3]~q ),
	.datad(!\sw_reset_ff_flush_counter[2]~q ),
	.datae(!\sw_reset_ff_flush~3_combout ),
	.dataf(!ff_rx_rdy),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush_counter[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush_counter[2]~2 .extended_lut = "off";
defparam \sw_reset_ff_flush_counter[2]~2 .lut_mask = 64'hFFFFFFFF7FFFFF7F;
defparam \sw_reset_ff_flush_counter[2]~2 .shared_arith = "off";

dffeas \sw_reset_ff_flush_counter[2] (
	.clk(clk_32_clk),
	.d(\sw_reset_ff_flush_counter[2]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sw_reset_ff_flush_counter[2]~q ),
	.prn(vcc));
defparam \sw_reset_ff_flush_counter[2] .is_wysiwyg = "true";
defparam \sw_reset_ff_flush_counter[2] .power_up = "low";

cyclonev_lcell_comb \sw_reset_ff_flush_counter[3]~1 (
	.dataa(!\sw_reset_ff_flush_counter[4]~q ),
	.datab(!\sw_reset_ff_flush~0_combout ),
	.datac(!\sw_reset_ff_flush_counter[3]~q ),
	.datad(!\sw_reset_ff_flush_counter[2]~q ),
	.datae(!\sw_reset_ff_flush~3_combout ),
	.dataf(!ff_rx_rdy),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush_counter[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush_counter[3]~1 .extended_lut = "off";
defparam \sw_reset_ff_flush_counter[3]~1 .lut_mask = 64'hFFFFFFFFF77F7FF7;
defparam \sw_reset_ff_flush_counter[3]~1 .shared_arith = "off";

dffeas \sw_reset_ff_flush_counter[3] (
	.clk(clk_32_clk),
	.d(\sw_reset_ff_flush_counter[3]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sw_reset_ff_flush_counter[3]~q ),
	.prn(vcc));
defparam \sw_reset_ff_flush_counter[3] .is_wysiwyg = "true";
defparam \sw_reset_ff_flush_counter[3] .power_up = "low";

cyclonev_lcell_comb \sw_reset_ff_flush~1 (
	.dataa(!\sw_reset_ff_flush_counter[3]~q ),
	.datab(!\sw_reset_ff_flush_counter[2]~q ),
	.datac(!\sw_reset_ff_flush_counter[1]~q ),
	.datad(!\sw_reset_ff_flush_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush~1 .extended_lut = "off";
defparam \sw_reset_ff_flush~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \sw_reset_ff_flush~1 .shared_arith = "off";

cyclonev_lcell_comb \sw_reset_ff_flush_counter[4]~0 (
	.dataa(!\sw_reset_ff_flush_counter[4]~q ),
	.datab(!\sw_reset_ff_flush~0_combout ),
	.datac(!\sw_reset_ff_flush~1_combout ),
	.datad(!ff_rx_rdy),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush_counter[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush_counter[4]~0 .extended_lut = "off";
defparam \sw_reset_ff_flush_counter[4]~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \sw_reset_ff_flush_counter[4]~0 .shared_arith = "off";

dffeas \sw_reset_ff_flush_counter[4] (
	.clk(clk_32_clk),
	.d(\sw_reset_ff_flush_counter[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sw_reset_ff_flush_counter[4]~q ),
	.prn(vcc));
defparam \sw_reset_ff_flush_counter[4] .is_wysiwyg = "true";
defparam \sw_reset_ff_flush_counter[4] .power_up = "low";

cyclonev_lcell_comb \sw_reset_ff_flush~2 (
	.dataa(!\sw_reset_ff_flush_counter[4]~q ),
	.datab(!\sw_reset_ff_flush~0_combout ),
	.datac(!\sw_reset_ff_flush~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sw_reset_ff_flush~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sw_reset_ff_flush~2 .extended_lut = "off";
defparam \sw_reset_ff_flush~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \sw_reset_ff_flush~2 .shared_arith = "off";

dffeas sw_reset_ff_flush(
	.clk(clk_32_clk),
	.d(\sw_reset_ff_flush~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sw_reset_ff_flush~q ),
	.prn(vcc));
defparam sw_reset_ff_flush.is_wysiwyg = "true";
defparam sw_reset_ff_flush.power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\Selector1~3_combout ),
	.datad(!\always10~0_combout ),
	.datae(!\state.LOC_STATE_WAIT~q ),
	.dataf(!\sw_reset_ff_flush~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hFFFFFFFFFFFBFFFF;
defparam \Selector2~0 .shared_arith = "off";

dffeas \state.LOC_STATE_WAIT (
	.clk(clk_32_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_WAIT~q ),
	.prn(vcc));
defparam \state.LOC_STATE_WAIT .is_wysiwyg = "true";
defparam \state.LOC_STATE_WAIT .power_up = "low";

cyclonev_lcell_comb \always10~1 (
	.dataa(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.datab(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.datac(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.datad(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.datae(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[21] ),
	.dataf(!\U_SYNC_5|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "off";
defparam \always10~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!sav_flag),
	.datac(!\rx_rdy_reg~q ),
	.datad(!\sw_reset_ff_flush~q ),
	.datae(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~0 .extended_lut = "off";
defparam \Selector0~0 .lut_mask = 64'hFFFFFFFFFFFFFFF6;
defparam \Selector0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!sav_flag),
	.datac(!\rx_rdy_reg~q ),
	.datad(!\state.LOC_STATE_WAIT~q ),
	.datae(!\sw_reset_ff_flush~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datac(!sav_flag),
	.datad(!\state.LOC_STATE_FF_DATA_FLUSH~q ),
	.datae(!\state.LOC_STATE_FF_DATA_FLUSH_WAIT~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \Selector9~0 .shared_arith = "off";

dffeas \state.LOC_STATE_FF_DATA_FLUSH_WAIT (
	.clk(clk_32_clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_FF_DATA_FLUSH_WAIT~q ),
	.prn(vcc));
defparam \state.LOC_STATE_FF_DATA_FLUSH_WAIT .is_wysiwyg = "true";
defparam \state.LOC_STATE_FF_DATA_FLUSH_WAIT .power_up = "low";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!\state.LOC_STATE_FF_DATA_FLUSH~q ),
	.datac(!\sw_reset_ff_flush~q ),
	.datad(!\state.LOC_STATE_IDLE~q ),
	.datae(!\state.LOC_STATE_FF_DATA_FLUSH_WAIT~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~2 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!sav_flag),
	.datac(!\state.LOC_STATE_IDLE~q ),
	.datad(!\always10~1_combout ),
	.datae(!\Selector5~0_combout ),
	.dataf(!\Selector5~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~2 .extended_lut = "off";
defparam \Selector5~2 .lut_mask = 64'hFFFFFFFFF7FFFFFF;
defparam \Selector5~2 .shared_arith = "off";

dffeas \state.LOC_STATE_FF_DATA_FLUSH (
	.clk(clk_32_clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_FF_DATA_FLUSH~q ),
	.prn(vcc));
defparam \state.LOC_STATE_FF_DATA_FLUSH .is_wysiwyg = "true";
defparam \state.LOC_STATE_FF_DATA_FLUSH .power_up = "low";

cyclonev_lcell_comb \Selector6~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!\state.LOC_STATE_FF_FLUSH_WAIT~q ),
	.datac(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datad(!\state.LOC_STATE_FF_DATA_FLUSH~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~0 .extended_lut = "off";
defparam \Selector6~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Selector6~0 .shared_arith = "off";

dffeas \state.LOC_STATE_FF_FLUSH_WAIT (
	.clk(clk_32_clk),
	.d(\Selector6~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_FF_FLUSH_WAIT~q ),
	.prn(vcc));
defparam \state.LOC_STATE_FF_FLUSH_WAIT .is_wysiwyg = "true";
defparam \state.LOC_STATE_FF_FLUSH_WAIT .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!stateLOC_STATE_SHIFT),
	.datab(!\RX_STATUS|empty_flag~q ),
	.datac(!\state.LOC_STATE_FF_FLUSH_WAIT~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Selector4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~2 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~2 .extended_lut = "off";
defparam \Selector4~2 .lut_mask = 64'hFFFFF7FFFFFFF7FF;
defparam \Selector4~2 .shared_arith = "off";

dffeas \state.LOC_STATE_END_FRM (
	.clk(clk_32_clk),
	.d(\Selector4~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_END_FRM~q ),
	.prn(vcc));
defparam \state.LOC_STATE_END_FRM .is_wysiwyg = "true";
defparam \state.LOC_STATE_END_FRM .power_up = "low";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!sav_flag),
	.datac(!\state.LOC_STATE_IDLE~q ),
	.datad(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\state.LOC_STATE_RST_DONE~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \Selector8~0 .shared_arith = "off";

dffeas \state.LOC_STATE_RST_DONE (
	.clk(clk_32_clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_RST_DONE~q ),
	.prn(vcc));
defparam \state.LOC_STATE_RST_DONE .is_wysiwyg = "true";
defparam \state.LOC_STATE_RST_DONE .power_up = "low";

cyclonev_lcell_comb \Selector0~1 (
	.dataa(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.datac(!\state.LOC_STATE_END_FRM~q ),
	.datad(!\state.LOC_STATE_RST_DONE~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~1 .extended_lut = "off";
defparam \Selector0~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \Selector0~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~2 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!\state.LOC_STATE_IDLE~q ),
	.datac(!\always10~1_combout ),
	.datad(!\Selector0~0_combout ),
	.datae(!\Selector0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~2 .extended_lut = "off";
defparam \Selector0~2 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \Selector0~2 .shared_arith = "off";

dffeas \state.LOC_STATE_IDLE (
	.clk(clk_32_clk),
	.d(\Selector0~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_IDLE~q ),
	.prn(vcc));
defparam \state.LOC_STATE_IDLE .is_wysiwyg = "true";
defparam \state.LOC_STATE_IDLE .power_up = "low";

cyclonev_lcell_comb \rx_err_sig~0 (
	.dataa(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.datab(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.datac(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.datad(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_err_sig~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_err_sig~0 .extended_lut = "off";
defparam \rx_err_sig~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \rx_err_sig~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!\RX_STATUS|empty_flag~q ),
	.datab(!\RX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[21] ),
	.datac(!\U_SYNC_5|std_sync_no_cut|dreg[1]~q ),
	.datad(!\state.LOC_STATE_IDLE~q ),
	.datae(!\rx_err_sig~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!\Selector1~0_combout ),
	.datab(!\always10~0_combout ),
	.datac(!\state.LOC_STATE_WAIT~q ),
	.datad(!\sw_reset_ff_flush~q ),
	.datae(!\Selector1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~0 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\rx_rdy_reg~q ),
	.dataf(!\state.LOC_STATE_SHIFT_WAIT~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~0 .extended_lut = "off";
defparam \Selector7~0 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \Selector7~0 .shared_arith = "off";

dffeas \state.LOC_STATE_SHIFT_WAIT (
	.clk(clk_32_clk),
	.d(\Selector7~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.LOC_STATE_SHIFT_WAIT~q ),
	.prn(vcc));
defparam \state.LOC_STATE_SHIFT_WAIT .is_wysiwyg = "true";
defparam \state.LOC_STATE_SHIFT_WAIT .power_up = "low";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\rx_rdy_reg~q ),
	.dataf(!\state.LOC_STATE_SHIFT_WAIT~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \rx_frm_type_reg~0 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_frm_type_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_frm_type_reg~0 .extended_lut = "off";
defparam \rx_frm_type_reg~0 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \rx_frm_type_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~1 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \Selector4~1 .shared_arith = "off";

cyclonev_lcell_comb \rx_frm_type_reg[1]~1 (
	.dataa(!stateLOC_STATE_SHIFT),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\Selector4~1_combout ),
	.datad(!\Selector4~0_combout ),
	.datae(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_frm_type_reg[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_frm_type_reg[1]~1 .extended_lut = "off";
defparam \rx_frm_type_reg[1]~1 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \rx_frm_type_reg[1]~1 .shared_arith = "off";

dffeas \rx_frm_type_reg[0] (
	.clk(clk_32_clk),
	.d(\rx_frm_type_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_frm_type_reg[1]~1_combout ),
	.q(\rx_frm_type_reg[0]~q ),
	.prn(vcc));
defparam \rx_frm_type_reg[0] .is_wysiwyg = "true";
defparam \rx_frm_type_reg[0] .power_up = "low";

cyclonev_lcell_comb \rx_frm_type_reg~2 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[36] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_frm_type_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_frm_type_reg~2 .extended_lut = "off";
defparam \rx_frm_type_reg~2 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \rx_frm_type_reg~2 .shared_arith = "off";

dffeas \rx_frm_type_reg[2] (
	.clk(clk_32_clk),
	.d(\rx_frm_type_reg~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_frm_type_reg[1]~1_combout ),
	.q(\rx_frm_type_reg[2]~q ),
	.prn(vcc));
defparam \rx_frm_type_reg[2] .is_wysiwyg = "true";
defparam \rx_frm_type_reg[2] .power_up = "low";

cyclonev_lcell_comb \rx_frm_type_reg~3 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_frm_type_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_frm_type_reg~3 .extended_lut = "off";
defparam \rx_frm_type_reg~3 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \rx_frm_type_reg~3 .shared_arith = "off";

dffeas \rx_frm_type_reg[1] (
	.clk(clk_32_clk),
	.d(\rx_frm_type_reg~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_frm_type_reg[1]~1_combout ),
	.q(\rx_frm_type_reg[1]~q ),
	.prn(vcc));
defparam \rx_frm_type_reg[1] .is_wysiwyg = "true";
defparam \rx_frm_type_reg[1] .power_up = "low";

cyclonev_lcell_comb \rx_frm_type_reg~4 (
	.dataa(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.datab(!stateLOC_STATE_DATA),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[39] ),
	.datae(!\Selector4~0_combout ),
	.dataf(!\RX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[37] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_frm_type_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_frm_type_reg~4 .extended_lut = "off";
defparam \rx_frm_type_reg~4 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \rx_frm_type_reg~4 .shared_arith = "off";

dffeas \rx_frm_type_reg[3] (
	.clk(clk_32_clk),
	.d(\rx_frm_type_reg~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rx_frm_type_reg[1]~1_combout ),
	.q(\rx_frm_type_reg[3]~q ),
	.prn(vcc));
defparam \rx_frm_type_reg[3] .is_wysiwyg = "true";
defparam \rx_frm_type_reg[3] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_35 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_35 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_35 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_36 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_36 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_36 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_37 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_37 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_37 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_38 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	rx_done_reg,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	rx_done_reg;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_38 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.rx_done_reg(rx_done_reg),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_38 (
	reset_n,
	dreg_1,
	rx_done_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	rx_done_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(!rx_done_reg),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_2 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_45 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_44 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_43 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_42 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_40 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_49 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_48 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_47 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_46 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_41 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_39 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_39 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_39 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_39 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_40 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_40 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_40 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_41 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_41 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_41 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_42 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_42 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_42 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_43 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_43 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_43 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_44 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_44 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_44 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_45 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_45 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_45 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_46 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_46 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_46 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_47 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_47 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_47 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_48 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_48 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_48 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_49 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_49 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_49 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_a_fifo_34 (
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_4,
	q_b_22,
	q_b_21,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	empty_flag1,
	Selector4,
	rx_stat_wren,
	payload_length_0,
	altera_tse_reset_synchronizer_chain_out,
	Selector41,
	payload_length_1,
	payload_length_2,
	payload_length_3,
	payload_length_4,
	payload_length_5,
	payload_length_6,
	payload_length_7,
	payload_length_8,
	payload_length_9,
	payload_length_10,
	payload_length_11,
	payload_length_12,
	payload_length_13,
	payload_length_14,
	payload_length_15,
	altera_tse_reset_synchronizer_chain_out1,
	Selector42,
	rx_stat_data_s_5,
	rx_stat_data_s_0,
	rx_stat_data_s_1,
	rx_stat_data_s_2,
	rx_stat_data_s_3,
	GND_port,
	clk_32_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_4;
output 	q_b_22;
output 	q_b_21;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	empty_flag1;
input 	Selector4;
input 	rx_stat_wren;
input 	payload_length_0;
input 	altera_tse_reset_synchronizer_chain_out;
input 	Selector41;
input 	payload_length_1;
input 	payload_length_2;
input 	payload_length_3;
input 	payload_length_4;
input 	payload_length_5;
input 	payload_length_6;
input 	payload_length_7;
input 	payload_length_8;
input 	payload_length_9;
input 	payload_length_10;
input 	payload_length_11;
input 	payload_length_12;
input 	payload_length_13;
input 	payload_length_14;
input 	payload_length_15;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	Selector42;
input 	rx_stat_data_s_5;
input 	rx_stat_data_s_0;
input 	rx_stat_data_s_1;
input 	rx_stat_data_s_2;
input 	rx_stat_data_s_3;
input 	GND_port;
input 	clk_32_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_WRT|b_out[0]~q ;
wire \U_WRT|b_out[1]~q ;
wire \U_WRT|b_out[2]~q ;
wire \U_WRT|b_out[3]~q ;
wire \U_WRT|b_out[4]~q ;
wire \U_WRT|b_out[5]~q ;
wire \U_WRT|b_out[6]~q ;
wire \U_WRT|b_out[7]~q ;
wire \U_WRT|b_out[8]~q ;
wire \U_RD|b_out[0]~q ;
wire \U_RD|b_out[1]~q ;
wire \U_RD|b_out[2]~q ;
wire \U_RD|b_out[3]~q ;
wire \U_RD|b_out[4]~q ;
wire \U_RD|b_out[5]~q ;
wire \U_RD|b_out[6]~q ;
wire \U_RD|b_out[7]~q ;
wire \U_RD|b_out[8]~q ;
wire \U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[5].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[6].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ;
wire \U_SYNC_WR_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ;
wire \wr_g_ptr_reg[4]~q ;
wire \wr_g_ptr_reg[5]~q ;
wire \wr_g_ptr_reg[6]~q ;
wire \wr_g_ptr_reg[7]~q ;
wire \wr_g_ptr_reg[8]~q ;
wire \wr_g_ptr_reg[1]~q ;
wire \wr_g_ptr_reg[2]~q ;
wire \wr_g_ptr_reg[3]~q ;
wire \wr_g_ptr_reg[0]~q ;
wire \U_WRT|g_out[4]~q ;
wire \U_WRT|g_out[5]~q ;
wire \U_WRT|g_out[6]~q ;
wire \U_WRT|g_out[7]~q ;
wire \U_WRT|g_out[8]~q ;
wire \U_WRT|g_out[1]~q ;
wire \U_WRT|g_out[2]~q ;
wire \U_WRT|g_out[3]~q ;
wire \U_WRT|g_out[0]~q ;
wire \ff_wr_binval[7]~3_combout ;
wire \wr_b_rptr[7]~q ;
wire \ff_wr_binval[5]~2_combout ;
wire \wr_b_rptr[6]~q ;
wire \ff_wr_binval[5]~1_combout ;
wire \wr_b_rptr[5]~q ;
wire \ff_wr_binval[3]~0_combout ;
wire \wr_b_rptr[4]~q ;
wire \ff_wr_binval[3]~4_combout ;
wire \wr_b_rptr[3]~q ;
wire \ff_wr_binval[1]~6_combout ;
wire \wr_b_rptr[2]~q ;
wire \ff_wr_binval[0]~5_combout ;
wire \wr_b_rptr[1]~q ;
wire \ff_wr_binval[0]~combout ;
wire \wr_b_rptr[0]~q ;
wire \ptr_rck_diff[0]~34 ;
wire \ptr_rck_diff[0]~35 ;
wire \ptr_rck_diff[1]~22 ;
wire \ptr_rck_diff[1]~23 ;
wire \ptr_rck_diff[2]~26 ;
wire \ptr_rck_diff[2]~27 ;
wire \ptr_rck_diff[3]~30 ;
wire \ptr_rck_diff[3]~31 ;
wire \ptr_rck_diff[4]~2 ;
wire \ptr_rck_diff[4]~3 ;
wire \ptr_rck_diff[5]~6 ;
wire \ptr_rck_diff[5]~7 ;
wire \ptr_rck_diff[6]~10 ;
wire \ptr_rck_diff[6]~11 ;
wire \ptr_rck_diff[7]~13_sumout ;
wire \wr_b_rptr[8]~q ;
wire \ptr_rck_diff[7]~14 ;
wire \ptr_rck_diff[7]~15 ;
wire \ptr_rck_diff[8]~17_sumout ;
wire \ptr_rck_diff[0]~33_sumout ;
wire \ptr_rck_diff[4]~1_sumout ;
wire \ptr_rck_diff[5]~5_sumout ;
wire \ptr_rck_diff[6]~9_sumout ;
wire \ptr_rck_diff[1]~21_sumout ;
wire \ptr_rck_diff[2]~25_sumout ;
wire \ptr_rck_diff[3]~29_sumout ;
wire \empty_flag~1_combout ;
wire \empty_flag~0_combout ;


IoTOctopus_QSYS_altera_tse_gray_cnt_2 U_WRT(
	.rx_stat_wren(rx_stat_wren),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo U_RAM(
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_16(q_b_16),
	.q_b_17(q_b_17),
	.q_b_18(q_b_18),
	.q_b_19(q_b_19),
	.q_b_20(q_b_20),
	.q_b_4(q_b_4),
	.q_b_22(q_b_22),
	.q_b_21(q_b_21),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.rx_stat_wren(rx_stat_wren),
	.payload_length_0(payload_length_0),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.b_out_01(\U_RD|b_out[0]~q ),
	.b_out_11(\U_RD|b_out[1]~q ),
	.b_out_21(\U_RD|b_out[2]~q ),
	.b_out_31(\U_RD|b_out[3]~q ),
	.b_out_41(\U_RD|b_out[4]~q ),
	.b_out_51(\U_RD|b_out[5]~q ),
	.b_out_61(\U_RD|b_out[6]~q ),
	.b_out_71(\U_RD|b_out[7]~q ),
	.b_out_81(\U_RD|b_out[8]~q ),
	.payload_length_1(payload_length_1),
	.payload_length_2(payload_length_2),
	.payload_length_3(payload_length_3),
	.payload_length_4(payload_length_4),
	.payload_length_5(payload_length_5),
	.payload_length_6(payload_length_6),
	.payload_length_7(payload_length_7),
	.payload_length_8(payload_length_8),
	.payload_length_9(payload_length_9),
	.payload_length_10(payload_length_10),
	.payload_length_11(payload_length_11),
	.payload_length_12(payload_length_12),
	.payload_length_13(payload_length_13),
	.payload_length_14(payload_length_14),
	.payload_length_15(payload_length_15),
	.rx_stat_data_s_5(rx_stat_data_s_5),
	.rx_stat_data_s_0(rx_stat_data_s_0),
	.rx_stat_data_s_1(rx_stat_data_s_1),
	.rx_stat_data_s_2(rx_stat_data_s_2),
	.rx_stat_data_s_3(rx_stat_data_s_3),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_4 U_SYNC_WR_G_PTR(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_01(\U_SYNC_WR_G_PTR|sync[5].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_02(\U_SYNC_WR_G_PTR|sync[6].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_03(\U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_04(\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_05(\U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_06(\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_07(\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.dreg_08(\U_SYNC_WR_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ),
	.wr_g_ptr_reg_4(\wr_g_ptr_reg[4]~q ),
	.wr_g_ptr_reg_5(\wr_g_ptr_reg[5]~q ),
	.wr_g_ptr_reg_6(\wr_g_ptr_reg[6]~q ),
	.wr_g_ptr_reg_7(\wr_g_ptr_reg[7]~q ),
	.wr_g_ptr_reg_8(\wr_g_ptr_reg[8]~q ),
	.wr_g_ptr_reg_1(\wr_g_ptr_reg[1]~q ),
	.wr_g_ptr_reg_2(\wr_g_ptr_reg[2]~q ),
	.wr_g_ptr_reg_3(\wr_g_ptr_reg[3]~q ),
	.wr_g_ptr_reg_0(\wr_g_ptr_reg[0]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_bin_cnt U_RD(
	.b_out_0(\U_RD|b_out[0]~q ),
	.b_out_1(\U_RD|b_out[1]~q ),
	.b_out_2(\U_RD|b_out[2]~q ),
	.b_out_3(\U_RD|b_out[3]~q ),
	.b_out_4(\U_RD|b_out[4]~q ),
	.b_out_5(\U_RD|b_out[5]~q ),
	.b_out_6(\U_RD|b_out[6]~q ),
	.b_out_7(\U_RD|b_out[7]~q ),
	.b_out_8(\U_RD|b_out[8]~q ),
	.reset(altera_tse_reset_synchronizer_chain_out),
	.clkena(Selector42),
	.clk(clk_32_clk));

dffeas \wr_g_ptr_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[4]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[4] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[4] .power_up = "low";

dffeas \wr_g_ptr_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[5]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[5] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[5] .power_up = "low";

dffeas \wr_g_ptr_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[6]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[6] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[6] .power_up = "low";

dffeas \wr_g_ptr_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[7]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[7] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[7] .power_up = "low";

dffeas \wr_g_ptr_reg[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[8]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[8] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[8] .power_up = "low";

dffeas \wr_g_ptr_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[1]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[1] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[1] .power_up = "low";

dffeas \wr_g_ptr_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[2]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[2] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[2] .power_up = "low";

dffeas \wr_g_ptr_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[3]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[3] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[3] .power_up = "low";

dffeas \wr_g_ptr_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_WRT|g_out[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_g_ptr_reg[0]~q ),
	.prn(vcc));
defparam \wr_g_ptr_reg[0] .is_wysiwyg = "true";
defparam \wr_g_ptr_reg[0] .power_up = "low";

dffeas empty_flag(
	.clk(clk_32_clk),
	.d(\empty_flag~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_flag1),
	.prn(vcc));
defparam empty_flag.is_wysiwyg = "true";
defparam empty_flag.power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[7]~3 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[7]~3 .extended_lut = "off";
defparam \ff_wr_binval[7]~3 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[7]~3 .shared_arith = "off";

dffeas \wr_b_rptr[7] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[7]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[7]~q ),
	.prn(vcc));
defparam \wr_b_rptr[7] .is_wysiwyg = "true";
defparam \wr_b_rptr[7] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[5]~2 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[6].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[5]~2 .extended_lut = "off";
defparam \ff_wr_binval[5]~2 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[5]~2 .shared_arith = "off";

dffeas \wr_b_rptr[6] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[6]~q ),
	.prn(vcc));
defparam \wr_b_rptr[6] .is_wysiwyg = "true";
defparam \wr_b_rptr[6] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[5]~1 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[5].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[6].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ),
	.datad(!\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[5]~1 .extended_lut = "off";
defparam \ff_wr_binval[5]~1 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[5]~1 .shared_arith = "off";

dffeas \wr_b_rptr[5] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[5]~q ),
	.prn(vcc));
defparam \wr_b_rptr[5] .is_wysiwyg = "true";
defparam \wr_b_rptr[5] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[3]~0 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[5].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[6].u|std_sync_no_cut|dreg[0]~q ),
	.datad(!\U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ),
	.datae(!\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~0 .extended_lut = "off";
defparam \ff_wr_binval[3]~0 .lut_mask = 64'h9669699696696996;
defparam \ff_wr_binval[3]~0 .shared_arith = "off";

dffeas \wr_b_rptr[4] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[4]~q ),
	.prn(vcc));
defparam \wr_b_rptr[4] .is_wysiwyg = "true";
defparam \wr_b_rptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[3]~4 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[3].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[4].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\U_SYNC_WR_G_PTR|sync[5].u|std_sync_no_cut|dreg[0]~q ),
	.datad(!\U_SYNC_WR_G_PTR|sync[6].u|std_sync_no_cut|dreg[0]~q ),
	.datae(!\U_SYNC_WR_G_PTR|sync[7].u|std_sync_no_cut|dreg[0]~q ),
	.dataf(!\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~4 .extended_lut = "off";
defparam \ff_wr_binval[3]~4 .lut_mask = 64'h6996966996696996;
defparam \ff_wr_binval[3]~4 .shared_arith = "off";

dffeas \wr_b_rptr[3] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[3]~q ),
	.prn(vcc));
defparam \wr_b_rptr[3] .is_wysiwyg = "true";
defparam \wr_b_rptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[1]~6 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\ff_wr_binval[3]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[1]~6 .extended_lut = "off";
defparam \ff_wr_binval[1]~6 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[1]~6 .shared_arith = "off";

dffeas \wr_b_rptr[2] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[1]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[2]~q ),
	.prn(vcc));
defparam \wr_b_rptr[2] .is_wysiwyg = "true";
defparam \wr_b_rptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0]~5 (
	.dataa(!\U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\ff_wr_binval[3]~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0]~5 .extended_lut = "off";
defparam \ff_wr_binval[0]~5 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[0]~5 .shared_arith = "off";

dffeas \wr_b_rptr[1] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[0]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[1]~q ),
	.prn(vcc));
defparam \wr_b_rptr[1] .is_wysiwyg = "true";
defparam \wr_b_rptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0] (
	.dataa(!\U_SYNC_WR_G_PTR|sync[1].u|std_sync_no_cut|dreg[0]~q ),
	.datab(!\U_SYNC_WR_G_PTR|sync[2].u|std_sync_no_cut|dreg[0]~q ),
	.datac(!\ff_wr_binval[3]~4_combout ),
	.datad(!\U_SYNC_WR_G_PTR|sync[0].u|std_sync_no_cut|dreg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0] .extended_lut = "off";
defparam \ff_wr_binval[0] .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[0] .shared_arith = "off";

dffeas \wr_b_rptr[0] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[0]~q ),
	.prn(vcc));
defparam \wr_b_rptr[0] .is_wysiwyg = "true";
defparam \wr_b_rptr[0] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[0]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[0]~q ),
	.datad(!\U_RD|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\ptr_rck_diff[0]~33_sumout ),
	.cout(\ptr_rck_diff[0]~34 ),
	.shareout(\ptr_rck_diff[0]~35 ));
defparam \ptr_rck_diff[0]~33 .extended_lut = "off";
defparam \ptr_rck_diff[0]~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[0]~33 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[1]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[1]~q ),
	.datad(!\U_RD|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[0]~34 ),
	.sharein(\ptr_rck_diff[0]~35 ),
	.combout(),
	.sumout(\ptr_rck_diff[1]~21_sumout ),
	.cout(\ptr_rck_diff[1]~22 ),
	.shareout(\ptr_rck_diff[1]~23 ));
defparam \ptr_rck_diff[1]~21 .extended_lut = "off";
defparam \ptr_rck_diff[1]~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[1]~21 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[2]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[2]~q ),
	.datad(!\U_RD|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[1]~22 ),
	.sharein(\ptr_rck_diff[1]~23 ),
	.combout(),
	.sumout(\ptr_rck_diff[2]~25_sumout ),
	.cout(\ptr_rck_diff[2]~26 ),
	.shareout(\ptr_rck_diff[2]~27 ));
defparam \ptr_rck_diff[2]~25 .extended_lut = "off";
defparam \ptr_rck_diff[2]~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[2]~25 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[3]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[3]~q ),
	.datad(!\U_RD|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[2]~26 ),
	.sharein(\ptr_rck_diff[2]~27 ),
	.combout(),
	.sumout(\ptr_rck_diff[3]~29_sumout ),
	.cout(\ptr_rck_diff[3]~30 ),
	.shareout(\ptr_rck_diff[3]~31 ));
defparam \ptr_rck_diff[3]~29 .extended_lut = "off";
defparam \ptr_rck_diff[3]~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[3]~29 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[4]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[4]~q ),
	.datad(!\U_RD|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[3]~30 ),
	.sharein(\ptr_rck_diff[3]~31 ),
	.combout(),
	.sumout(\ptr_rck_diff[4]~1_sumout ),
	.cout(\ptr_rck_diff[4]~2 ),
	.shareout(\ptr_rck_diff[4]~3 ));
defparam \ptr_rck_diff[4]~1 .extended_lut = "off";
defparam \ptr_rck_diff[4]~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[4]~1 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[5]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[5]~q ),
	.datad(!\U_RD|b_out[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[4]~2 ),
	.sharein(\ptr_rck_diff[4]~3 ),
	.combout(),
	.sumout(\ptr_rck_diff[5]~5_sumout ),
	.cout(\ptr_rck_diff[5]~6 ),
	.shareout(\ptr_rck_diff[5]~7 ));
defparam \ptr_rck_diff[5]~5 .extended_lut = "off";
defparam \ptr_rck_diff[5]~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[5]~5 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[6]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[6]~q ),
	.datad(!\U_RD|b_out[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[5]~6 ),
	.sharein(\ptr_rck_diff[5]~7 ),
	.combout(),
	.sumout(\ptr_rck_diff[6]~9_sumout ),
	.cout(\ptr_rck_diff[6]~10 ),
	.shareout(\ptr_rck_diff[6]~11 ));
defparam \ptr_rck_diff[6]~9 .extended_lut = "off";
defparam \ptr_rck_diff[6]~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[6]~9 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[7]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[7]~q ),
	.datad(!\U_RD|b_out[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[6]~10 ),
	.sharein(\ptr_rck_diff[6]~11 ),
	.combout(),
	.sumout(\ptr_rck_diff[7]~13_sumout ),
	.cout(\ptr_rck_diff[7]~14 ),
	.shareout(\ptr_rck_diff[7]~15 ));
defparam \ptr_rck_diff[7]~13 .extended_lut = "off";
defparam \ptr_rck_diff[7]~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[7]~13 .shared_arith = "on";

dffeas \wr_b_rptr[8] (
	.clk(clk_32_clk),
	.d(\U_SYNC_WR_G_PTR|sync[8].u|std_sync_no_cut|dreg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[8]~q ),
	.prn(vcc));
defparam \wr_b_rptr[8] .is_wysiwyg = "true";
defparam \wr_b_rptr[8] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[8]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[8]~q ),
	.datad(!\U_RD|b_out[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[7]~14 ),
	.sharein(\ptr_rck_diff[7]~15 ),
	.combout(),
	.sumout(\ptr_rck_diff[8]~17_sumout ),
	.cout(),
	.shareout());
defparam \ptr_rck_diff[8]~17 .extended_lut = "off";
defparam \ptr_rck_diff[8]~17 .lut_mask = 64'h0000000000000FF0;
defparam \ptr_rck_diff[8]~17 .shared_arith = "on";

cyclonev_lcell_comb \empty_flag~1 (
	.dataa(!\ptr_rck_diff[4]~1_sumout ),
	.datab(!\ptr_rck_diff[5]~5_sumout ),
	.datac(!\ptr_rck_diff[6]~9_sumout ),
	.datad(!\ptr_rck_diff[1]~21_sumout ),
	.datae(!\ptr_rck_diff[2]~25_sumout ),
	.dataf(!\ptr_rck_diff[3]~29_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~1 .extended_lut = "off";
defparam \empty_flag~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \empty_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \empty_flag~0 (
	.dataa(!\ptr_rck_diff[7]~13_sumout ),
	.datab(!\ptr_rck_diff[8]~17_sumout ),
	.datac(!Selector41),
	.datad(!Selector4),
	.datae(!\ptr_rck_diff[0]~33_sumout ),
	.dataf(!\empty_flag~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~0 .extended_lut = "off";
defparam \empty_flag~0 .lut_mask = 64'hFFFFFFFFF7FFFFFF;
defparam \empty_flag~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_4 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	dreg_01,
	dreg_02,
	dreg_03,
	dreg_04,
	dreg_05,
	dreg_06,
	dreg_07,
	dreg_08,
	wr_g_ptr_reg_4,
	wr_g_ptr_reg_5,
	wr_g_ptr_reg_6,
	wr_g_ptr_reg_7,
	wr_g_ptr_reg_8,
	wr_g_ptr_reg_1,
	wr_g_ptr_reg_2,
	wr_g_ptr_reg_3,
	wr_g_ptr_reg_0,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
output 	dreg_01;
output 	dreg_02;
output 	dreg_03;
output 	dreg_04;
output 	dreg_05;
output 	dreg_06;
output 	dreg_07;
output 	dreg_08;
input 	wr_g_ptr_reg_4;
input 	wr_g_ptr_reg_5;
input 	wr_g_ptr_reg_6;
input 	wr_g_ptr_reg_7;
input 	wr_g_ptr_reg_8;
input 	wr_g_ptr_reg_1;
input 	wr_g_ptr_reg_2;
input 	wr_g_ptr_reg_3;
input 	wr_g_ptr_reg_0;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_69 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_04),
	.wr_g_ptr_reg_8(wr_g_ptr_reg_8),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_68 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_03),
	.wr_g_ptr_reg_7(wr_g_ptr_reg_7),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_67 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_02),
	.wr_g_ptr_reg_6(wr_g_ptr_reg_6),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_66 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_01),
	.wr_g_ptr_reg_5(wr_g_ptr_reg_5),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_65 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.wr_g_ptr_reg_4(wr_g_ptr_reg_4),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_64 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_07),
	.wr_g_ptr_reg_3(wr_g_ptr_reg_3),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_63 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_06),
	.wr_g_ptr_reg_2(wr_g_ptr_reg_2),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_62 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_05),
	.wr_g_ptr_reg_1(wr_g_ptr_reg_1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_61 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_08),
	.wr_g_ptr_reg_0(wr_g_ptr_reg_0),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_61 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_0,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_0;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_61 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_0),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_61 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_62 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_62 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_62 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_63 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_2,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_2;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_63 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_2),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_63 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_64 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_3,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_3;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_64 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_3),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_64 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_65 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_4,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_4;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_65 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_4),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_65 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_66 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_5,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_5;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_66 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_5),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_66 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_67 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_6,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_6;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_67 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_6),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_67 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_68 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_7,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_7;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_68 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_7),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_68 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_69 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_0,
	wr_g_ptr_reg_8,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_0;
input 	wr_g_ptr_reg_8;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_69 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_0(dreg_0),
	.din(wr_g_ptr_reg_8),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_69 (
	reset_n,
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo (
	q_b_5,
	q_b_6,
	q_b_7,
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_16,
	q_b_17,
	q_b_18,
	q_b_19,
	q_b_20,
	q_b_4,
	q_b_22,
	q_b_21,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	rx_stat_wren,
	payload_length_0,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	b_out_01,
	b_out_11,
	b_out_21,
	b_out_31,
	b_out_41,
	b_out_51,
	b_out_61,
	b_out_71,
	b_out_81,
	payload_length_1,
	payload_length_2,
	payload_length_3,
	payload_length_4,
	payload_length_5,
	payload_length_6,
	payload_length_7,
	payload_length_8,
	payload_length_9,
	payload_length_10,
	payload_length_11,
	payload_length_12,
	payload_length_13,
	payload_length_14,
	payload_length_15,
	rx_stat_data_s_5,
	rx_stat_data_s_0,
	rx_stat_data_s_1,
	rx_stat_data_s_2,
	rx_stat_data_s_3,
	GND_port,
	clk_32_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_16;
output 	q_b_17;
output 	q_b_18;
output 	q_b_19;
output 	q_b_20;
output 	q_b_4;
output 	q_b_22;
output 	q_b_21;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
input 	rx_stat_wren;
input 	payload_length_0;
input 	b_out_0;
input 	b_out_1;
input 	b_out_2;
input 	b_out_3;
input 	b_out_4;
input 	b_out_5;
input 	b_out_6;
input 	b_out_7;
input 	b_out_8;
input 	b_out_01;
input 	b_out_11;
input 	b_out_21;
input 	b_out_31;
input 	b_out_41;
input 	b_out_51;
input 	b_out_61;
input 	b_out_71;
input 	b_out_81;
input 	payload_length_1;
input 	payload_length_2;
input 	payload_length_3;
input 	payload_length_4;
input 	payload_length_5;
input 	payload_length_6;
input 	payload_length_7;
input 	payload_length_8;
input 	payload_length_9;
input 	payload_length_10;
input 	payload_length_11;
input 	payload_length_12;
input 	payload_length_13;
input 	payload_length_14;
input 	payload_length_15;
input 	rx_stat_data_s_5;
input 	rx_stat_data_s_0;
input 	rx_stat_data_s_1;
input 	rx_stat_data_s_2;
input 	rx_stat_data_s_3;
input 	GND_port;
input 	clk_32_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_2 altsyncram_component(
	.q_b({q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_unconnected_wire_35,q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,
q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,
q_b_1,q_b_0}),
	.wren_a(rx_stat_wren),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,GND_port,rx_stat_data_s_5,payload_length_15,payload_length_14,payload_length_13,payload_length_12,payload_length_11,payload_length_10,payload_length_9,payload_length_8,payload_length_7,payload_length_6,
payload_length_5,payload_length_4,payload_length_3,payload_length_2,payload_length_1,payload_length_0,gnd,rx_stat_data_s_3,rx_stat_data_s_2,rx_stat_data_s_1,rx_stat_data_s_0}),
	.address_a({gnd,gnd,b_out_8,b_out_7,b_out_6,b_out_5,b_out_4,b_out_3,b_out_2,b_out_1,b_out_0}),
	.address_b({gnd,gnd,b_out_81,b_out_71,b_out_61,b_out_51,b_out_41,b_out_31,b_out_21,b_out_11,b_out_01}),
	.clock1(clk_32_clk),
	.clock0(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altsyncram_2 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	wren_a;
input 	[39:0] data_a;
input 	[10:0] address_a;
input 	[10:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_t3o1 auto_generated(
	.q_b({q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[22],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock1(clock1),
	.clock0(clock0));

endmodule

module IoTOctopus_QSYS_altsyncram_t3o1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[22:0] q_b;
input 	wren_a;
input 	[22:0] data_a;
input 	[8:0] address_a;
input 	[8:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 9;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 511;
defparam ram_block1a5.port_a_logical_ram_depth = 512;
defparam ram_block1a5.port_a_logical_ram_width = 23;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 9;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 511;
defparam ram_block1a5.port_b_logical_ram_depth = 512;
defparam ram_block1a5.port_b_logical_ram_width = 23;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 9;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 511;
defparam ram_block1a6.port_a_logical_ram_depth = 512;
defparam ram_block1a6.port_a_logical_ram_width = 23;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 9;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 511;
defparam ram_block1a6.port_b_logical_ram_depth = 512;
defparam ram_block1a6.port_b_logical_ram_width = 23;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 9;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 511;
defparam ram_block1a7.port_a_logical_ram_depth = 512;
defparam ram_block1a7.port_a_logical_ram_width = 23;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 9;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 511;
defparam ram_block1a7.port_b_logical_ram_depth = 512;
defparam ram_block1a7.port_b_logical_ram_width = 23;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 9;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 511;
defparam ram_block1a8.port_a_logical_ram_depth = 512;
defparam ram_block1a8.port_a_logical_ram_width = 23;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 9;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 511;
defparam ram_block1a8.port_b_logical_ram_depth = 512;
defparam ram_block1a8.port_b_logical_ram_width = 23;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 9;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 511;
defparam ram_block1a9.port_a_logical_ram_depth = 512;
defparam ram_block1a9.port_a_logical_ram_width = 23;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 9;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 511;
defparam ram_block1a9.port_b_logical_ram_depth = 512;
defparam ram_block1a9.port_b_logical_ram_width = 23;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 9;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 511;
defparam ram_block1a10.port_a_logical_ram_depth = 512;
defparam ram_block1a10.port_a_logical_ram_width = 23;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 9;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 511;
defparam ram_block1a10.port_b_logical_ram_depth = 512;
defparam ram_block1a10.port_b_logical_ram_width = 23;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 9;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 511;
defparam ram_block1a11.port_a_logical_ram_depth = 512;
defparam ram_block1a11.port_a_logical_ram_width = 23;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 9;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 511;
defparam ram_block1a11.port_b_logical_ram_depth = 512;
defparam ram_block1a11.port_b_logical_ram_width = 23;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 9;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 511;
defparam ram_block1a12.port_a_logical_ram_depth = 512;
defparam ram_block1a12.port_a_logical_ram_width = 23;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 9;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 511;
defparam ram_block1a12.port_b_logical_ram_depth = 512;
defparam ram_block1a12.port_b_logical_ram_width = 23;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 9;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 511;
defparam ram_block1a13.port_a_logical_ram_depth = 512;
defparam ram_block1a13.port_a_logical_ram_width = 23;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 9;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 511;
defparam ram_block1a13.port_b_logical_ram_depth = 512;
defparam ram_block1a13.port_b_logical_ram_width = 23;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 9;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 511;
defparam ram_block1a14.port_a_logical_ram_depth = 512;
defparam ram_block1a14.port_a_logical_ram_width = 23;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 9;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 511;
defparam ram_block1a14.port_b_logical_ram_depth = 512;
defparam ram_block1a14.port_b_logical_ram_width = 23;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 9;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 511;
defparam ram_block1a15.port_a_logical_ram_depth = 512;
defparam ram_block1a15.port_a_logical_ram_width = 23;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 9;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 511;
defparam ram_block1a15.port_b_logical_ram_depth = 512;
defparam ram_block1a15.port_b_logical_ram_width = 23;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 9;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 511;
defparam ram_block1a16.port_a_logical_ram_depth = 512;
defparam ram_block1a16.port_a_logical_ram_width = 23;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 9;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 511;
defparam ram_block1a16.port_b_logical_ram_depth = 512;
defparam ram_block1a16.port_b_logical_ram_width = 23;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 9;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 511;
defparam ram_block1a17.port_a_logical_ram_depth = 512;
defparam ram_block1a17.port_a_logical_ram_width = 23;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 9;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 511;
defparam ram_block1a17.port_b_logical_ram_depth = 512;
defparam ram_block1a17.port_b_logical_ram_width = 23;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 9;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 511;
defparam ram_block1a18.port_a_logical_ram_depth = 512;
defparam ram_block1a18.port_a_logical_ram_width = 23;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 9;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 511;
defparam ram_block1a18.port_b_logical_ram_depth = 512;
defparam ram_block1a18.port_b_logical_ram_width = 23;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 9;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 511;
defparam ram_block1a19.port_a_logical_ram_depth = 512;
defparam ram_block1a19.port_a_logical_ram_width = 23;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 9;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 511;
defparam ram_block1a19.port_b_logical_ram_depth = 512;
defparam ram_block1a19.port_b_logical_ram_width = 23;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 9;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 511;
defparam ram_block1a20.port_a_logical_ram_depth = 512;
defparam ram_block1a20.port_a_logical_ram_width = 23;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 9;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 511;
defparam ram_block1a20.port_b_logical_ram_depth = 512;
defparam ram_block1a20.port_b_logical_ram_width = 23;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 9;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 511;
defparam ram_block1a4.port_a_logical_ram_depth = 512;
defparam ram_block1a4.port_a_logical_ram_width = 23;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 9;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 511;
defparam ram_block1a4.port_b_logical_ram_depth = 512;
defparam ram_block1a4.port_b_logical_ram_width = 23;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 9;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 511;
defparam ram_block1a22.port_a_logical_ram_depth = 512;
defparam ram_block1a22.port_a_logical_ram_width = 23;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 9;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 511;
defparam ram_block1a22.port_b_logical_ram_depth = 512;
defparam ram_block1a22.port_b_logical_ram_width = 23;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 9;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 511;
defparam ram_block1a21.port_a_logical_ram_depth = 512;
defparam ram_block1a21.port_a_logical_ram_width = 23;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 9;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 511;
defparam ram_block1a21.port_b_logical_ram_depth = 512;
defparam ram_block1a21.port_b_logical_ram_width = 23;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 9;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 511;
defparam ram_block1a0.port_a_logical_ram_depth = 512;
defparam ram_block1a0.port_a_logical_ram_width = 23;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 9;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 511;
defparam ram_block1a0.port_b_logical_ram_depth = 512;
defparam ram_block1a0.port_b_logical_ram_width = 23;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 9;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 511;
defparam ram_block1a1.port_a_logical_ram_depth = 512;
defparam ram_block1a1.port_a_logical_ram_width = 23;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 9;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 511;
defparam ram_block1a1.port_b_logical_ram_depth = 512;
defparam ram_block1a1.port_b_logical_ram_width = 23;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 9;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 511;
defparam ram_block1a2.port_a_logical_ram_depth = 512;
defparam ram_block1a2.port_a_logical_ram_width = 23;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 9;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 511;
defparam ram_block1a2.port_b_logical_ram_depth = 512;
defparam ram_block1a2.port_b_logical_ram_width = 23;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_34:RX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_t3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 9;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 511;
defparam ram_block1a3.port_a_logical_ram_depth = 512;
defparam ram_block1a3.port_a_logical_ram_width = 23;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 9;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 511;
defparam ram_block1a3.port_b_logical_ram_depth = 512;
defparam ram_block1a3.port_b_logical_ram_width = 23;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module IoTOctopus_QSYS_altera_tse_bin_cnt (
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	reset,
	clkena,
	clk)/* synthesis synthesis_greybox=1 */;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	b_out_5;
output 	b_out_6;
output 	b_out_7;
output 	b_out_8;
input 	reset;
input 	clkena;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \b_int[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \b_int[3]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \b_int[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \b_int[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \b_int[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \b_int[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \b_int[8]~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \b_int[1]~q ;
wire \Add0~1_sumout ;
wire \b_int~0_combout ;
wire \b_int[0]~q ;
wire \b_out[0]~0_combout ;


dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[5] (
	.clk(clk),
	.d(\b_int[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[6] (
	.clk(clk),
	.d(\b_int[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[7] (
	.clk(clk),
	.d(\b_int[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \b_int[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \b_int[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[5]~q ),
	.prn(vcc));
defparam \b_int[5] .is_wysiwyg = "true";
defparam \b_int[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \b_int[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[6]~q ),
	.prn(vcc));
defparam \b_int[6] .is_wysiwyg = "true";
defparam \b_int[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \b_int[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[7]~q ),
	.prn(vcc));
defparam \b_int[7] .is_wysiwyg = "true";
defparam \b_int[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \b_int[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[8]~q ),
	.prn(vcc));
defparam \b_int[8] .is_wysiwyg = "true";
defparam \b_int[8] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[4]~q ),
	.datac(!\b_int[5]~q ),
	.datad(!\b_int[6]~q ),
	.datae(!\b_int[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(!\b_int[3]~q ),
	.datad(!\b_int[8]~q ),
	.datae(!\LessThan0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan0~1 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \b_int~0 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(!\b_int[3]~q ),
	.datad(!\b_int[8]~q ),
	.datae(!\Add0~1_sumout ),
	.dataf(!\LessThan0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int~0 .extended_lut = "off";
defparam \b_int~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \b_int~0 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clkena),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_2 (
	rx_stat_wren,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	reset,
	g_out_4,
	g_out_5,
	g_out_6,
	g_out_7,
	g_out_8,
	g_out_1,
	g_out_2,
	g_out_3,
	g_out_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rx_stat_wren;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	b_out_5;
output 	b_out_6;
output 	b_out_7;
output 	b_out_8;
input 	reset;
output 	g_out_4;
output 	g_out_5;
output 	g_out_6;
output 	g_out_7;
output 	g_out_8;
output 	g_out_1;
output 	g_out_2;
output 	g_out_3;
output 	g_out_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \b_int[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \b_int[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \b_int[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \b_int[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \b_int[8]~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \b_int[1]~q ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \b_int[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \b_int[3]~q ;
wire \Add0~1_sumout ;
wire \b_int~0_combout ;
wire \b_int[0]~q ;
wire \b_out[0]~0_combout ;
wire \gry_grayval[4]~combout ;
wire \gry_grayval[5]~combout ;
wire \gry_grayval[6]~combout ;
wire \gry_grayval[7]~combout ;
wire \gry_grayval[1]~combout ;
wire \gry_grayval[2]~combout ;
wire \gry_grayval[3]~combout ;
wire \gry_grayval[0]~combout ;


dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[5] (
	.clk(clk),
	.d(\b_int[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[6] (
	.clk(clk),
	.d(\b_int[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[7] (
	.clk(clk),
	.d(\b_int[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

dffeas \g_out[4] (
	.clk(clk),
	.d(\gry_grayval[4]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[5] (
	.clk(clk),
	.d(\gry_grayval[5]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_5),
	.prn(vcc));
defparam \g_out[5] .is_wysiwyg = "true";
defparam \g_out[5] .power_up = "low";

dffeas \g_out[6] (
	.clk(clk),
	.d(\gry_grayval[6]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_6),
	.prn(vcc));
defparam \g_out[6] .is_wysiwyg = "true";
defparam \g_out[6] .power_up = "low";

dffeas \g_out[7] (
	.clk(clk),
	.d(\gry_grayval[7]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_7),
	.prn(vcc));
defparam \g_out[7] .is_wysiwyg = "true";
defparam \g_out[7] .power_up = "low";

dffeas \g_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_8),
	.prn(vcc));
defparam \g_out[8] .is_wysiwyg = "true";
defparam \g_out[8] .power_up = "low";

dffeas \g_out[1] (
	.clk(clk),
	.d(\gry_grayval[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[2] (
	.clk(clk),
	.d(\gry_grayval[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[3] (
	.clk(clk),
	.d(\gry_grayval[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[0] (
	.clk(clk),
	.d(\gry_grayval[0]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \b_int[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[5]~q ),
	.prn(vcc));
defparam \b_int[5] .is_wysiwyg = "true";
defparam \b_int[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \b_int[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[6]~q ),
	.prn(vcc));
defparam \b_int[6] .is_wysiwyg = "true";
defparam \b_int[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \b_int[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[7]~q ),
	.prn(vcc));
defparam \b_int[7] .is_wysiwyg = "true";
defparam \b_int[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \b_int[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[8]~q ),
	.prn(vcc));
defparam \b_int[8] .is_wysiwyg = "true";
defparam \b_int[8] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(!\b_int[2]~q ),
	.datad(!\b_int[6]~q ),
	.datae(!\b_int[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(!\b_int[5]~q ),
	.datad(!\b_int[7]~q ),
	.datae(!\LessThan0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan0~1 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

dffeas \b_int[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \b_int~0 (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(!\b_int[5]~q ),
	.datad(!\b_int[7]~q ),
	.datae(!\Add0~1_sumout ),
	.dataf(!\LessThan0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int~0 .extended_lut = "off";
defparam \b_int~0 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \b_int~0 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_stat_wren),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[4] (
	.dataa(!\b_int[4]~q ),
	.datab(!\b_int[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[4] .extended_lut = "off";
defparam \gry_grayval[4] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[4] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[5] (
	.dataa(!\b_int[5]~q ),
	.datab(!\b_int[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[5] .extended_lut = "off";
defparam \gry_grayval[5] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[5] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[6] (
	.dataa(!\b_int[6]~q ),
	.datab(!\b_int[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[6] .extended_lut = "off";
defparam \gry_grayval[6] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[6] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[7] (
	.dataa(!\b_int[7]~q ),
	.datab(!\b_int[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[7] .extended_lut = "off";
defparam \gry_grayval[7] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[7] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[1] (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[1] .extended_lut = "off";
defparam \gry_grayval[1] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[1] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[2] (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[2] .extended_lut = "off";
defparam \gry_grayval[2] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[2] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[3] (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[3] .extended_lut = "off";
defparam \gry_grayval[3] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[3] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[0] (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[0] .extended_lut = "off";
defparam \gry_grayval[0] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[0] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_a_fifo_opt_1246 (
	q_b_32,
	q_b_39,
	q_b_34,
	q_b_33,
	q_b_36,
	q_b_35,
	q_b_37,
	sav_flag1,
	afull_flag1,
	aempty_flag1,
	rx_wren32,
	rx_eop32,
	altera_tse_reset_synchronizer_chain_out,
	byte_empty_1,
	frm_type32_0,
	rx_sop32,
	frm_type32_2,
	frm_type32_1,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	altera_tse_reset_synchronizer_chain_out1,
	data_rdreq,
	GND_port,
	clk_32_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_32;
output 	q_b_39;
output 	q_b_34;
output 	q_b_33;
output 	q_b_36;
output 	q_b_35;
output 	q_b_37;
output 	sav_flag1;
output 	afull_flag1;
output 	aempty_flag1;
input 	rx_wren32;
input 	rx_eop32;
input 	altera_tse_reset_synchronizer_chain_out;
input 	byte_empty_1;
input 	frm_type32_0;
input 	rx_sop32;
input 	frm_type32_2;
input 	frm_type32_1;
input 	dreg_1;
input 	dreg_11;
input 	dreg_12;
input 	dreg_13;
input 	dreg_14;
input 	dreg_15;
input 	dreg_16;
input 	dreg_17;
input 	dreg_18;
input 	dreg_19;
input 	dreg_110;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	data_rdreq;
input 	GND_port;
input 	clk_32_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_WRT|b_out[0]~q ;
wire \U_WRT|b_out[1]~q ;
wire \U_WRT|b_out[2]~q ;
wire \U_WRT|b_out[3]~q ;
wire \U_WRT|b_out[4]~q ;
wire \U_WRT|b_out[5]~q ;
wire \U_WRT|b_out[6]~q ;
wire \U_WRT|b_out[7]~q ;
wire \U_WRT|b_out[8]~q ;
wire \U_WRT|b_out[9]~q ;
wire \U_WRT|b_out[10]~q ;
wire \U_RD|b_out[0]~q ;
wire \U_RD|b_out[1]~q ;
wire \U_RD|b_out[2]~q ;
wire \U_RD|b_out[3]~q ;
wire \U_RD|b_out[4]~q ;
wire \U_RD|b_out[5]~q ;
wire \U_RD|b_out[6]~q ;
wire \U_RD|b_out[7]~q ;
wire \U_RD|b_out[8]~q ;
wire \U_RD|b_out[9]~q ;
wire \U_RD|b_out[10]~q ;
wire \U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_WRT|g_out[10]~q ;
wire \U_WRT|g_out[9]~q ;
wire \U_WRT|g_out[8]~q ;
wire \U_WRT|g_out[7]~q ;
wire \U_WRT|g_out[6]~q ;
wire \U_WRT|g_out[5]~q ;
wire \U_WRT|g_out[4]~q ;
wire \U_WRT|g_out[3]~q ;
wire \U_WRT|g_out[2]~q ;
wire \U_WRT|g_out[1]~q ;
wire \U_WRT|g_out[0]~q ;
wire \U_RD|g_out[10]~q ;
wire \U_RD|g_out[9]~q ;
wire \U_RD|g_out[8]~q ;
wire \U_RD|g_out[7]~q ;
wire \U_RD|g_out[6]~q ;
wire \U_RD|g_out[5]~q ;
wire \U_RD|g_out[4]~q ;
wire \U_RD|g_out[3]~q ;
wire \U_RD|g_out[2]~q ;
wire \U_RD|g_out[0]~q ;
wire \U_RD|g_out[1]~q ;
wire \wr_b_rptr[10]~q ;
wire \ff_wr_binval[9]~7_combout ;
wire \wr_b_rptr[9]~q ;
wire \ff_wr_binval[8]~8_combout ;
wire \wr_b_rptr[8]~q ;
wire \ff_wr_binval[6]~5_combout ;
wire \wr_b_rptr[7]~q ;
wire \ff_wr_binval[6]~6_combout ;
wire \wr_b_rptr[6]~q ;
wire \ff_wr_binval[4]~0_combout ;
wire \wr_b_rptr[5]~q ;
wire \ff_wr_binval[4]~4_combout ;
wire \wr_b_rptr[4]~q ;
wire \ff_wr_binval[3]~2_combout ;
wire \wr_b_rptr[3]~q ;
wire \ff_wr_binval[1]~3_combout ;
wire \wr_b_rptr[2]~q ;
wire \ff_wr_binval[0]~1_combout ;
wire \wr_b_rptr[1]~q ;
wire \ff_wr_binval[0]~combout ;
wire \wr_b_rptr[0]~q ;
wire \Add1~10 ;
wire \Add1~11 ;
wire \Add1~6 ;
wire \Add1~7 ;
wire \Add1~18 ;
wire \Add1~19 ;
wire \Add1~14 ;
wire \Add1~15 ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~22 ;
wire \Add1~23 ;
wire \Add1~34 ;
wire \Add1~35 ;
wire \Add1~30 ;
wire \Add1~31 ;
wire \Add1~42 ;
wire \Add1~43 ;
wire \Add1~38 ;
wire \Add1~39 ;
wire \Add1~1_sumout ;
wire \ptr_rck_diff[10]~q ;
wire \LessThan4~0_combout ;
wire \Add1~5_sumout ;
wire \ptr_rck_diff[1]~q ;
wire \Add1~9_sumout ;
wire \ptr_rck_diff[0]~q ;
wire \LessThan4~1_combout ;
wire \Add1~13_sumout ;
wire \ptr_rck_diff[3]~q ;
wire \Add1~17_sumout ;
wire \ptr_rck_diff[2]~q ;
wire \LessThan4~2_combout ;
wire \LessThan4~3_combout ;
wire \Add1~21_sumout ;
wire \ptr_rck_diff[5]~q ;
wire \Add1~25_sumout ;
wire \ptr_rck_diff[4]~q ;
wire \LessThan4~4_combout ;
wire \LessThan4~5_combout ;
wire \Add1~29_sumout ;
wire \ptr_rck_diff[7]~q ;
wire \Add1~33_sumout ;
wire \ptr_rck_diff[6]~q ;
wire \LessThan4~6_combout ;
wire \LessThan4~7_combout ;
wire \LessThan4~8_combout ;
wire \Add1~37_sumout ;
wire \ptr_rck_diff[9]~q ;
wire \Add1~41_sumout ;
wire \ptr_rck_diff[8]~q ;
wire \sav_flag~0_combout ;
wire \sav_flag~1_combout ;
wire \Equal5~0_combout ;
wire \Equal5~1_combout ;
wire \sav_flag~2_combout ;
wire \sav_flag~3_combout ;
wire \rd_b_wptr[10]~q ;
wire \ff_rd_binval[9]~7_combout ;
wire \rd_b_wptr[9]~q ;
wire \ff_rd_binval[8]~8_combout ;
wire \rd_b_wptr[8]~q ;
wire \ff_rd_binval[6]~5_combout ;
wire \rd_b_wptr[7]~q ;
wire \ff_rd_binval[6]~6_combout ;
wire \rd_b_wptr[6]~q ;
wire \ff_rd_binval[4]~0_combout ;
wire \rd_b_wptr[5]~q ;
wire \ff_rd_binval[4]~4_combout ;
wire \rd_b_wptr[4]~q ;
wire \ff_rd_binval[3]~2_combout ;
wire \rd_b_wptr[3]~q ;
wire \ff_rd_binval[1]~3_combout ;
wire \rd_b_wptr[2]~q ;
wire \ff_rd_binval[0]~1_combout ;
wire \rd_b_wptr[1]~q ;
wire \ff_rd_binval[0]~combout ;
wire \rd_b_wptr[0]~q ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~1_sumout ;
wire \ptr_wck_diff[10]~q ;
wire \LessThan0~0_combout ;
wire \Add0~5_sumout ;
wire \ptr_wck_diff[0]~q ;
wire \Add0~9_sumout ;
wire \ptr_wck_diff[1]~q ;
wire \LessThan0~1_combout ;
wire \Add0~13_sumout ;
wire \ptr_wck_diff[3]~q ;
wire \Add0~17_sumout ;
wire \ptr_wck_diff[2]~q ;
wire \LessThan0~2_combout ;
wire \LessThan0~3_combout ;
wire \Add0~21_sumout ;
wire \ptr_wck_diff[5]~q ;
wire \Add0~25_sumout ;
wire \ptr_wck_diff[4]~q ;
wire \LessThan0~4_combout ;
wire \LessThan0~5_combout ;
wire \Add0~29_sumout ;
wire \ptr_wck_diff[7]~q ;
wire \Add0~33_sumout ;
wire \ptr_wck_diff[6]~q ;
wire \LessThan0~6_combout ;
wire \LessThan0~7_combout ;
wire \LessThan0~8_combout ;
wire \Add0~37_sumout ;
wire \ptr_wck_diff[9]~q ;
wire \Add0~41_sumout ;
wire \ptr_wck_diff[8]~q ;
wire \afull_flag~0_combout ;
wire \afull_flag~1_combout ;
wire \afull_flag~2_combout ;
wire \afull_flag~3_combout ;
wire \afull_flag~4_combout ;
wire \afull_flag~5_combout ;
wire \LessThan3~0_combout ;
wire \LessThan3~1_combout ;
wire \LessThan3~2_combout ;
wire \LessThan3~3_combout ;
wire \LessThan3~4_combout ;
wire \LessThan3~5_combout ;
wire \LessThan3~6_combout ;
wire \LessThan3~7_combout ;
wire \LessThan3~8_combout ;
wire \aempty_flag~0_combout ;
wire \aempty_flag~1_combout ;
wire \aempty_flag~2_combout ;
wire \aempty_flag~3_combout ;
wire \aempty_flag~4_combout ;
wire \aempty_flag~5_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_8 U_SYNC_4(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_7 U_SYNC_3(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_3|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.g_out_10(\U_WRT|g_out[10]~q ),
	.g_out_9(\U_WRT|g_out[9]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_6 U_SYNC_2(
	.dreg_1(\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_5 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.g_out_10(\U_RD|g_out[10]~q ),
	.g_out_9(\U_RD|g_out[9]~q ),
	.g_out_8(\U_RD|g_out[8]~q ),
	.g_out_7(\U_RD|g_out[7]~q ),
	.g_out_6(\U_RD|g_out[6]~q ),
	.g_out_5(\U_RD|g_out[5]~q ),
	.g_out_4(\U_RD|g_out[4]~q ),
	.g_out_3(\U_RD|g_out[3]~q ),
	.g_out_2(\U_RD|g_out[2]~q ),
	.g_out_0(\U_RD|g_out[0]~q ),
	.g_out_1(\U_RD|g_out[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_3 U_RD(
	.b_out_0(\U_RD|b_out[0]~q ),
	.b_out_1(\U_RD|b_out[1]~q ),
	.b_out_2(\U_RD|b_out[2]~q ),
	.b_out_3(\U_RD|b_out[3]~q ),
	.b_out_4(\U_RD|b_out[4]~q ),
	.b_out_5(\U_RD|b_out[5]~q ),
	.b_out_6(\U_RD|b_out[6]~q ),
	.b_out_7(\U_RD|b_out[7]~q ),
	.b_out_8(\U_RD|b_out[8]~q ),
	.b_out_9(\U_RD|b_out[9]~q ),
	.b_out_10(\U_RD|b_out[10]~q ),
	.reset(altera_tse_reset_synchronizer_chain_out),
	.data_rdreq(data_rdreq),
	.g_out_10(\U_RD|g_out[10]~q ),
	.g_out_9(\U_RD|g_out[9]~q ),
	.g_out_8(\U_RD|g_out[8]~q ),
	.g_out_7(\U_RD|g_out[7]~q ),
	.g_out_6(\U_RD|g_out[6]~q ),
	.g_out_5(\U_RD|g_out[5]~q ),
	.g_out_4(\U_RD|g_out[4]~q ),
	.g_out_3(\U_RD|g_out[3]~q ),
	.g_out_2(\U_RD|g_out[2]~q ),
	.g_out_0(\U_RD|g_out[0]~q ),
	.g_out_1(\U_RD|g_out[1]~q ),
	.clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_4 U_WRT(
	.rx_wren32(rx_wren32),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.b_out_9(\U_WRT|b_out[9]~q ),
	.b_out_10(\U_WRT|b_out[10]~q ),
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.g_out_10(\U_WRT|g_out[10]~q ),
	.g_out_9(\U_WRT|g_out[9]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_1 U_RAM(
	.q_b_32(q_b_32),
	.q_b_39(q_b_39),
	.q_b_34(q_b_34),
	.q_b_33(q_b_33),
	.q_b_36(q_b_36),
	.q_b_35(q_b_35),
	.q_b_37(q_b_37),
	.rx_wren32(rx_wren32),
	.rx_eop32(rx_eop32),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.b_out_9(\U_WRT|b_out[9]~q ),
	.b_out_10(\U_WRT|b_out[10]~q ),
	.b_out_01(\U_RD|b_out[0]~q ),
	.b_out_11(\U_RD|b_out[1]~q ),
	.b_out_21(\U_RD|b_out[2]~q ),
	.b_out_31(\U_RD|b_out[3]~q ),
	.b_out_41(\U_RD|b_out[4]~q ),
	.b_out_51(\U_RD|b_out[5]~q ),
	.b_out_61(\U_RD|b_out[6]~q ),
	.b_out_71(\U_RD|b_out[7]~q ),
	.b_out_81(\U_RD|b_out[8]~q ),
	.b_out_91(\U_RD|b_out[9]~q ),
	.b_out_101(\U_RD|b_out[10]~q ),
	.byte_empty_1(byte_empty_1),
	.frm_type32_0(frm_type32_0),
	.rx_sop32(rx_sop32),
	.frm_type32_2(frm_type32_2),
	.frm_type32_1(frm_type32_1),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

dffeas sav_flag(
	.clk(clk_32_clk),
	.d(\sav_flag~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sav_flag1),
	.prn(vcc));
defparam sav_flag.is_wysiwyg = "true";
defparam sav_flag.power_up = "low";

dffeas afull_flag(
	.clk(mac_rx_clock_connection_clk),
	.d(\afull_flag~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(afull_flag1),
	.prn(vcc));
defparam afull_flag.is_wysiwyg = "true";
defparam afull_flag.power_up = "low";

dffeas aempty_flag(
	.clk(clk_32_clk),
	.d(\aempty_flag~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(aempty_flag1),
	.prn(vcc));
defparam aempty_flag.is_wysiwyg = "true";
defparam aempty_flag.power_up = "low";

dffeas \wr_b_rptr[10] (
	.clk(clk_32_clk),
	.d(\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[10]~q ),
	.prn(vcc));
defparam \wr_b_rptr[10] .is_wysiwyg = "true";
defparam \wr_b_rptr[10] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[9]~7 (
	.dataa(!\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[9]~7 .extended_lut = "off";
defparam \ff_wr_binval[9]~7 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[9]~7 .shared_arith = "off";

dffeas \wr_b_rptr[9] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[9]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[9]~q ),
	.prn(vcc));
defparam \wr_b_rptr[9] .is_wysiwyg = "true";
defparam \wr_b_rptr[9] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[8]~8 (
	.dataa(!\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[8]~8 .extended_lut = "off";
defparam \ff_wr_binval[8]~8 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[8]~8 .shared_arith = "off";

dffeas \wr_b_rptr[8] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[8]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[8]~q ),
	.prn(vcc));
defparam \wr_b_rptr[8] .is_wysiwyg = "true";
defparam \wr_b_rptr[8] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[6]~5 (
	.dataa(!\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[6]~5 .extended_lut = "off";
defparam \ff_wr_binval[6]~5 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[6]~5 .shared_arith = "off";

dffeas \wr_b_rptr[7] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[7]~q ),
	.prn(vcc));
defparam \wr_b_rptr[7] .is_wysiwyg = "true";
defparam \wr_b_rptr[7] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[6]~6 (
	.dataa(!\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[6]~6 .extended_lut = "off";
defparam \ff_wr_binval[6]~6 .lut_mask = 64'h9669699696696996;
defparam \ff_wr_binval[6]~6 .shared_arith = "off";

dffeas \wr_b_rptr[6] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[6]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[6]~q ),
	.prn(vcc));
defparam \wr_b_rptr[6] .is_wysiwyg = "true";
defparam \wr_b_rptr[6] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[4]~0 (
	.dataa(!\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_3|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[4]~0 .extended_lut = "off";
defparam \ff_wr_binval[4]~0 .lut_mask = 64'h6996966996696996;
defparam \ff_wr_binval[4]~0 .shared_arith = "off";

dffeas \wr_b_rptr[5] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[5]~q ),
	.prn(vcc));
defparam \wr_b_rptr[5] .is_wysiwyg = "true";
defparam \wr_b_rptr[5] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[4]~4 (
	.dataa(!\ff_wr_binval[4]~0_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[4]~4 .extended_lut = "off";
defparam \ff_wr_binval[4]~4 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[4]~4 .shared_arith = "off";

dffeas \wr_b_rptr[4] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[4]~q ),
	.prn(vcc));
defparam \wr_b_rptr[4] .is_wysiwyg = "true";
defparam \wr_b_rptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[3]~2 (
	.dataa(!\ff_wr_binval[4]~0_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~2 .extended_lut = "off";
defparam \ff_wr_binval[3]~2 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[3]~2 .shared_arith = "off";

dffeas \wr_b_rptr[3] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[3]~q ),
	.prn(vcc));
defparam \wr_b_rptr[3] .is_wysiwyg = "true";
defparam \wr_b_rptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[1]~3 (
	.dataa(!\ff_wr_binval[4]~0_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[1]~3 .extended_lut = "off";
defparam \ff_wr_binval[1]~3 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[1]~3 .shared_arith = "off";

dffeas \wr_b_rptr[2] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[2]~q ),
	.prn(vcc));
defparam \wr_b_rptr[2] .is_wysiwyg = "true";
defparam \wr_b_rptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0]~1 (
	.dataa(!\ff_wr_binval[4]~0_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0]~1 .extended_lut = "off";
defparam \ff_wr_binval[0]~1 .lut_mask = 64'h9669699696696996;
defparam \ff_wr_binval[0]~1 .shared_arith = "off";

dffeas \wr_b_rptr[1] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[1]~q ),
	.prn(vcc));
defparam \wr_b_rptr[1] .is_wysiwyg = "true";
defparam \wr_b_rptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0] (
	.dataa(!\ff_wr_binval[4]~0_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0] .extended_lut = "off";
defparam \ff_wr_binval[0] .lut_mask = 64'h6996966996696996;
defparam \ff_wr_binval[0] .shared_arith = "off";

dffeas \wr_b_rptr[0] (
	.clk(clk_32_clk),
	.d(\ff_wr_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[0]~q ),
	.prn(vcc));
defparam \wr_b_rptr[0] .is_wysiwyg = "true";
defparam \wr_b_rptr[0] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[0]~q ),
	.datad(!\U_RD|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout(\Add1~11 ));
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~9 .shared_arith = "on";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[1]~q ),
	.datad(!\U_RD|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(\Add1~11 ),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout(\Add1~7 ));
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~5 .shared_arith = "on";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[2]~q ),
	.datad(!\U_RD|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(\Add1~7 ),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout(\Add1~19 ));
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~17 .shared_arith = "on";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[3]~q ),
	.datad(!\U_RD|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(\Add1~19 ),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout(\Add1~15 ));
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~13 .shared_arith = "on";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[4]~q ),
	.datad(!\U_RD|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(\Add1~15 ),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout(\Add1~27 ));
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~25 .shared_arith = "on";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[5]~q ),
	.datad(!\U_RD|b_out[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(\Add1~27 ),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout(\Add1~23 ));
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~21 .shared_arith = "on";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[6]~q ),
	.datad(!\U_RD|b_out[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(\Add1~23 ),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout(\Add1~35 ));
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~33 .shared_arith = "on";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[7]~q ),
	.datad(!\U_RD|b_out[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(\Add1~35 ),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout(\Add1~31 ));
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~29 .shared_arith = "on";

cyclonev_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[8]~q ),
	.datad(!\U_RD|b_out[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(\Add1~31 ),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout(\Add1~43 ));
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~41 .shared_arith = "on";

cyclonev_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[9]~q ),
	.datad(!\U_RD|b_out[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(\Add1~43 ),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout(\Add1~39 ));
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~37 .shared_arith = "on";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[10]~q ),
	.datad(!\U_RD|b_out[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(\Add1~39 ),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000000000000FF0;
defparam \Add1~1 .shared_arith = "on";

dffeas \ptr_rck_diff[10] (
	.clk(clk_32_clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[10]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[10] .is_wysiwyg = "true";
defparam \ptr_rck_diff[10] .power_up = "low";

cyclonev_lcell_comb \LessThan4~0 (
	.dataa(!dreg_1),
	.datab(!\ptr_rck_diff[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~0 .extended_lut = "off";
defparam \LessThan4~0 .lut_mask = 64'h6666666666666666;
defparam \LessThan4~0 .shared_arith = "off";

dffeas \ptr_rck_diff[1] (
	.clk(clk_32_clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[1]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[1] .is_wysiwyg = "true";
defparam \ptr_rck_diff[1] .power_up = "low";

dffeas \ptr_rck_diff[0] (
	.clk(clk_32_clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[0]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[0] .is_wysiwyg = "true";
defparam \ptr_rck_diff[0] .power_up = "low";

cyclonev_lcell_comb \LessThan4~1 (
	.dataa(!dreg_11),
	.datab(!dreg_12),
	.datac(!\ptr_rck_diff[1]~q ),
	.datad(!\ptr_rck_diff[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~1 .extended_lut = "off";
defparam \LessThan4~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan4~1 .shared_arith = "off";

dffeas \ptr_rck_diff[3] (
	.clk(clk_32_clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[3]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[3] .is_wysiwyg = "true";
defparam \ptr_rck_diff[3] .power_up = "low";

dffeas \ptr_rck_diff[2] (
	.clk(clk_32_clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[2]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[2] .is_wysiwyg = "true";
defparam \ptr_rck_diff[2] .power_up = "low";

cyclonev_lcell_comb \LessThan4~2 (
	.dataa(!dreg_13),
	.datab(!dreg_14),
	.datac(!\ptr_rck_diff[3]~q ),
	.datad(!\ptr_rck_diff[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~2 .extended_lut = "off";
defparam \LessThan4~2 .lut_mask = 64'h6996699669966996;
defparam \LessThan4~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~3 (
	.dataa(!dreg_13),
	.datab(!dreg_14),
	.datac(!\ptr_rck_diff[3]~q ),
	.datad(!\ptr_rck_diff[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~3 .extended_lut = "off";
defparam \LessThan4~3 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan4~3 .shared_arith = "off";

dffeas \ptr_rck_diff[5] (
	.clk(clk_32_clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[5]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[5] .is_wysiwyg = "true";
defparam \ptr_rck_diff[5] .power_up = "low";

dffeas \ptr_rck_diff[4] (
	.clk(clk_32_clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[4]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[4] .is_wysiwyg = "true";
defparam \ptr_rck_diff[4] .power_up = "low";

cyclonev_lcell_comb \LessThan4~4 (
	.dataa(!dreg_15),
	.datab(!dreg_16),
	.datac(!\ptr_rck_diff[5]~q ),
	.datad(!\ptr_rck_diff[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~4 .extended_lut = "off";
defparam \LessThan4~4 .lut_mask = 64'h6996699669966996;
defparam \LessThan4~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~5 (
	.dataa(!dreg_15),
	.datab(!dreg_16),
	.datac(!\ptr_rck_diff[5]~q ),
	.datad(!\ptr_rck_diff[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~5 .extended_lut = "off";
defparam \LessThan4~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan4~5 .shared_arith = "off";

dffeas \ptr_rck_diff[7] (
	.clk(clk_32_clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[7]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[7] .is_wysiwyg = "true";
defparam \ptr_rck_diff[7] .power_up = "low";

dffeas \ptr_rck_diff[6] (
	.clk(clk_32_clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[6]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[6] .is_wysiwyg = "true";
defparam \ptr_rck_diff[6] .power_up = "low";

cyclonev_lcell_comb \LessThan4~6 (
	.dataa(!dreg_17),
	.datab(!dreg_18),
	.datac(!\ptr_rck_diff[7]~q ),
	.datad(!\ptr_rck_diff[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~6 .extended_lut = "off";
defparam \LessThan4~6 .lut_mask = 64'h6996699669966996;
defparam \LessThan4~6 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~7 (
	.dataa(!\LessThan4~1_combout ),
	.datab(!\LessThan4~2_combout ),
	.datac(!\LessThan4~3_combout ),
	.datad(!\LessThan4~4_combout ),
	.datae(!\LessThan4~5_combout ),
	.dataf(!\LessThan4~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~7 .extended_lut = "off";
defparam \LessThan4~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \LessThan4~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~8 (
	.dataa(!dreg_17),
	.datab(!dreg_18),
	.datac(!\ptr_rck_diff[7]~q ),
	.datad(!\ptr_rck_diff[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~8 .extended_lut = "off";
defparam \LessThan4~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan4~8 .shared_arith = "off";

dffeas \ptr_rck_diff[9] (
	.clk(clk_32_clk),
	.d(\Add1~37_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[9]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[9] .is_wysiwyg = "true";
defparam \ptr_rck_diff[9] .power_up = "low";

dffeas \ptr_rck_diff[8] (
	.clk(clk_32_clk),
	.d(\Add1~41_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[8]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[8] .is_wysiwyg = "true";
defparam \ptr_rck_diff[8] .power_up = "low";

cyclonev_lcell_comb \sav_flag~0 (
	.dataa(!dreg_19),
	.datab(!dreg_110),
	.datac(!\ptr_rck_diff[9]~q ),
	.datad(!\ptr_rck_diff[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~0 .extended_lut = "off";
defparam \sav_flag~0 .lut_mask = 64'h6996699669966996;
defparam \sav_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \sav_flag~1 (
	.dataa(!dreg_19),
	.datab(!dreg_110),
	.datac(!\ptr_rck_diff[9]~q ),
	.datad(!\ptr_rck_diff[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~1 .extended_lut = "off";
defparam \sav_flag~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sav_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!dreg_11),
	.datab(!dreg_12),
	.datac(!dreg_13),
	.datad(!dreg_14),
	.datae(!dreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~1 (
	.dataa(!dreg_17),
	.datab(!dreg_18),
	.datac(!dreg_19),
	.datad(!dreg_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~1 .extended_lut = "off";
defparam \Equal5~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal5~1 .shared_arith = "off";

cyclonev_lcell_comb \sav_flag~2 (
	.dataa(!dreg_16),
	.datab(!dreg_1),
	.datac(!\ptr_rck_diff[10]~q ),
	.datad(!\Equal5~0_combout ),
	.datae(!\Equal5~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~2 .extended_lut = "off";
defparam \sav_flag~2 .lut_mask = 64'hB8FFFFFFB8FFFFFF;
defparam \sav_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \sav_flag~3 (
	.dataa(!\LessThan4~0_combout ),
	.datab(!\LessThan4~7_combout ),
	.datac(!\LessThan4~8_combout ),
	.datad(!\sav_flag~0_combout ),
	.datae(!\sav_flag~1_combout ),
	.dataf(!\sav_flag~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~3 .extended_lut = "off";
defparam \sav_flag~3 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \sav_flag~3 .shared_arith = "off";

dffeas \rd_b_wptr[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[10]~q ),
	.prn(vcc));
defparam \rd_b_wptr[10] .is_wysiwyg = "true";
defparam \rd_b_wptr[10] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[9]~7 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[9]~7 .extended_lut = "off";
defparam \ff_rd_binval[9]~7 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[9]~7 .shared_arith = "off";

dffeas \rd_b_wptr[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[9]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[9]~q ),
	.prn(vcc));
defparam \rd_b_wptr[9] .is_wysiwyg = "true";
defparam \rd_b_wptr[9] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[8]~8 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[8]~8 .extended_lut = "off";
defparam \ff_rd_binval[8]~8 .lut_mask = 64'h9696969696969696;
defparam \ff_rd_binval[8]~8 .shared_arith = "off";

dffeas \rd_b_wptr[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[8]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[8]~q ),
	.prn(vcc));
defparam \rd_b_wptr[8] .is_wysiwyg = "true";
defparam \rd_b_wptr[8] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[6]~5 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[6]~5 .extended_lut = "off";
defparam \ff_rd_binval[6]~5 .lut_mask = 64'h6996699669966996;
defparam \ff_rd_binval[6]~5 .shared_arith = "off";

dffeas \rd_b_wptr[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[7]~q ),
	.prn(vcc));
defparam \rd_b_wptr[7] .is_wysiwyg = "true";
defparam \rd_b_wptr[7] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[6]~6 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[6]~6 .extended_lut = "off";
defparam \ff_rd_binval[6]~6 .lut_mask = 64'h9669699696696996;
defparam \ff_rd_binval[6]~6 .shared_arith = "off";

dffeas \rd_b_wptr[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[6]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[6]~q ),
	.prn(vcc));
defparam \rd_b_wptr[6] .is_wysiwyg = "true";
defparam \rd_b_wptr[6] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[4]~0 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[4]~0 .extended_lut = "off";
defparam \ff_rd_binval[4]~0 .lut_mask = 64'h6996966996696996;
defparam \ff_rd_binval[4]~0 .shared_arith = "off";

dffeas \rd_b_wptr[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[5]~q ),
	.prn(vcc));
defparam \rd_b_wptr[5] .is_wysiwyg = "true";
defparam \rd_b_wptr[5] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[4]~4 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[4]~4 .extended_lut = "off";
defparam \ff_rd_binval[4]~4 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[4]~4 .shared_arith = "off";

dffeas \rd_b_wptr[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[4]~q ),
	.prn(vcc));
defparam \rd_b_wptr[4] .is_wysiwyg = "true";
defparam \rd_b_wptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[3]~2 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[3]~2 .extended_lut = "off";
defparam \ff_rd_binval[3]~2 .lut_mask = 64'h9696969696969696;
defparam \ff_rd_binval[3]~2 .shared_arith = "off";

dffeas \rd_b_wptr[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[3]~q ),
	.prn(vcc));
defparam \rd_b_wptr[3] .is_wysiwyg = "true";
defparam \rd_b_wptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[1]~3 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[1]~3 .extended_lut = "off";
defparam \ff_rd_binval[1]~3 .lut_mask = 64'h6996699669966996;
defparam \ff_rd_binval[1]~3 .shared_arith = "off";

dffeas \rd_b_wptr[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[2]~q ),
	.prn(vcc));
defparam \rd_b_wptr[2] .is_wysiwyg = "true";
defparam \rd_b_wptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[0]~1 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[0]~1 .extended_lut = "off";
defparam \ff_rd_binval[0]~1 .lut_mask = 64'h9669699696696996;
defparam \ff_rd_binval[0]~1 .shared_arith = "off";

dffeas \rd_b_wptr[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[1]~q ),
	.prn(vcc));
defparam \rd_b_wptr[1] .is_wysiwyg = "true";
defparam \rd_b_wptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[0] (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[0] .extended_lut = "off";
defparam \ff_rd_binval[0] .lut_mask = 64'h6996966996696996;
defparam \ff_rd_binval[0] .shared_arith = "off";

dffeas \rd_b_wptr[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ff_rd_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[0]~q ),
	.prn(vcc));
defparam \rd_b_wptr[0] .is_wysiwyg = "true";
defparam \rd_b_wptr[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[0]~q ),
	.datad(!\U_WRT|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[1]~q ),
	.datad(!\U_WRT|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[2]~q ),
	.datad(!\U_WRT|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[3]~q ),
	.datad(!\U_WRT|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[4]~q ),
	.datad(!\U_WRT|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[5]~q ),
	.datad(!\U_WRT|b_out[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[6]~q ),
	.datad(!\U_WRT|b_out[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[7]~q ),
	.datad(!\U_WRT|b_out[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[8]~q ),
	.datad(!\U_WRT|b_out[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[9]~q ),
	.datad(!\U_WRT|b_out[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[10]~q ),
	.datad(!\U_WRT|b_out[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000000000000FF0;
defparam \Add0~1 .shared_arith = "on";

dffeas \ptr_wck_diff[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[10]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[10] .is_wysiwyg = "true";
defparam \ptr_wck_diff[10] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\ptr_wck_diff[10]~q ),
	.datab(!\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h6666666666666666;
defparam \LessThan0~0 .shared_arith = "off";

dffeas \ptr_wck_diff[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[0]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[0] .is_wysiwyg = "true";
defparam \ptr_wck_diff[0] .power_up = "low";

dffeas \ptr_wck_diff[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[1]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[1] .is_wysiwyg = "true";
defparam \ptr_wck_diff[1] .power_up = "low";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\ptr_wck_diff[0]~q ),
	.datab(!\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[1]~q ),
	.datad(!\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

dffeas \ptr_wck_diff[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[3]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[3] .is_wysiwyg = "true";
defparam \ptr_wck_diff[3] .power_up = "low";

dffeas \ptr_wck_diff[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[2]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[2] .is_wysiwyg = "true";
defparam \ptr_wck_diff[2] .power_up = "low";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!\ptr_wck_diff[3]~q ),
	.datab(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[2]~q ),
	.datad(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h6996699669966996;
defparam \LessThan0~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~3 (
	.dataa(!\ptr_wck_diff[3]~q ),
	.datab(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[2]~q ),
	.datad(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~3 .extended_lut = "off";
defparam \LessThan0~3 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~3 .shared_arith = "off";

dffeas \ptr_wck_diff[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[5]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[5] .is_wysiwyg = "true";
defparam \ptr_wck_diff[5] .power_up = "low";

dffeas \ptr_wck_diff[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[4]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[4] .is_wysiwyg = "true";
defparam \ptr_wck_diff[4] .power_up = "low";

cyclonev_lcell_comb \LessThan0~4 (
	.dataa(!\ptr_wck_diff[5]~q ),
	.datab(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[4]~q ),
	.datad(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~4 .extended_lut = "off";
defparam \LessThan0~4 .lut_mask = 64'h6996699669966996;
defparam \LessThan0~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~5 (
	.dataa(!\ptr_wck_diff[5]~q ),
	.datab(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[4]~q ),
	.datad(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~5 .extended_lut = "off";
defparam \LessThan0~5 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~5 .shared_arith = "off";

dffeas \ptr_wck_diff[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[7]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[7] .is_wysiwyg = "true";
defparam \ptr_wck_diff[7] .power_up = "low";

dffeas \ptr_wck_diff[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[6]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[6] .is_wysiwyg = "true";
defparam \ptr_wck_diff[6] .power_up = "low";

cyclonev_lcell_comb \LessThan0~6 (
	.dataa(!\ptr_wck_diff[7]~q ),
	.datab(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[6]~q ),
	.datad(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~6 .extended_lut = "off";
defparam \LessThan0~6 .lut_mask = 64'h6996699669966996;
defparam \LessThan0~6 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~7 (
	.dataa(!\LessThan0~1_combout ),
	.datab(!\LessThan0~2_combout ),
	.datac(!\LessThan0~3_combout ),
	.datad(!\LessThan0~4_combout ),
	.datae(!\LessThan0~5_combout ),
	.dataf(!\LessThan0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~7 .extended_lut = "off";
defparam \LessThan0~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \LessThan0~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~8 (
	.dataa(!\ptr_wck_diff[7]~q ),
	.datab(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[6]~q ),
	.datad(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~8 .extended_lut = "off";
defparam \LessThan0~8 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~8 .shared_arith = "off";

dffeas \ptr_wck_diff[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[9]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[9] .is_wysiwyg = "true";
defparam \ptr_wck_diff[9] .power_up = "low";

dffeas \ptr_wck_diff[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[8]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[8] .is_wysiwyg = "true";
defparam \ptr_wck_diff[8] .power_up = "low";

cyclonev_lcell_comb \afull_flag~0 (
	.dataa(!\ptr_wck_diff[9]~q ),
	.datab(!\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[8]~q ),
	.datad(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~0 .extended_lut = "off";
defparam \afull_flag~0 .lut_mask = 64'h6996699669966996;
defparam \afull_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~1 (
	.dataa(!\ptr_wck_diff[9]~q ),
	.datab(!\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_wck_diff[8]~q ),
	.datad(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~1 .extended_lut = "off";
defparam \afull_flag~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \afull_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~2 (
	.dataa(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~2 .extended_lut = "off";
defparam \afull_flag~2 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \afull_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~3 (
	.dataa(!\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~3 .extended_lut = "off";
defparam \afull_flag~3 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \afull_flag~3 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~4 (
	.dataa(!\ptr_wck_diff[10]~q ),
	.datab(!\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\afull_flag~2_combout ),
	.datae(!\afull_flag~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~4 .extended_lut = "off";
defparam \afull_flag~4 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \afull_flag~4 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~5 (
	.dataa(!\LessThan0~0_combout ),
	.datab(!\LessThan0~7_combout ),
	.datac(!\LessThan0~8_combout ),
	.datad(!\afull_flag~0_combout ),
	.datae(!\afull_flag~1_combout ),
	.dataf(!\afull_flag~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~5 .extended_lut = "off";
defparam \afull_flag~5 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \afull_flag~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!\ptr_rck_diff[10]~q ),
	.datab(!\U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h6666666666666666;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~1 (
	.dataa(!\ptr_rck_diff[1]~q ),
	.datab(!\ptr_rck_diff[0]~q ),
	.datac(!\U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~1 .extended_lut = "off";
defparam \LessThan3~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan3~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~2 (
	.dataa(!\ptr_rck_diff[3]~q ),
	.datab(!\ptr_rck_diff[2]~q ),
	.datac(!\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~2 .extended_lut = "off";
defparam \LessThan3~2 .lut_mask = 64'h6996699669966996;
defparam \LessThan3~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~3 (
	.dataa(!\ptr_rck_diff[3]~q ),
	.datab(!\ptr_rck_diff[2]~q ),
	.datac(!\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~3 .extended_lut = "off";
defparam \LessThan3~3 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan3~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~4 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\ptr_rck_diff[4]~q ),
	.datac(!\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~4 .extended_lut = "off";
defparam \LessThan3~4 .lut_mask = 64'h6996699669966996;
defparam \LessThan3~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~5 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\ptr_rck_diff[4]~q ),
	.datac(!\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~5 .extended_lut = "off";
defparam \LessThan3~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan3~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~6 (
	.dataa(!\ptr_rck_diff[7]~q ),
	.datab(!\ptr_rck_diff[6]~q ),
	.datac(!\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~6 .extended_lut = "off";
defparam \LessThan3~6 .lut_mask = 64'h6996699669966996;
defparam \LessThan3~6 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~7 (
	.dataa(!\LessThan3~1_combout ),
	.datab(!\LessThan3~2_combout ),
	.datac(!\LessThan3~3_combout ),
	.datad(!\LessThan3~4_combout ),
	.datae(!\LessThan3~5_combout ),
	.dataf(!\LessThan3~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~7 .extended_lut = "off";
defparam \LessThan3~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \LessThan3~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~8 (
	.dataa(!\ptr_rck_diff[7]~q ),
	.datab(!\ptr_rck_diff[6]~q ),
	.datac(!\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~8 .extended_lut = "off";
defparam \LessThan3~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan3~8 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~0 (
	.dataa(!\ptr_rck_diff[9]~q ),
	.datab(!\ptr_rck_diff[8]~q ),
	.datac(!\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~0 .extended_lut = "off";
defparam \aempty_flag~0 .lut_mask = 64'h6996699669966996;
defparam \aempty_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~1 (
	.dataa(!\ptr_rck_diff[9]~q ),
	.datab(!\ptr_rck_diff[8]~q ),
	.datac(!\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~1 .extended_lut = "off";
defparam \aempty_flag~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \aempty_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~2 (
	.dataa(!\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~2 .extended_lut = "off";
defparam \aempty_flag~2 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \aempty_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~3 (
	.dataa(!\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~3 .extended_lut = "off";
defparam \aempty_flag~3 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \aempty_flag~3 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~4 (
	.dataa(!\ptr_rck_diff[10]~q ),
	.datab(!\U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\aempty_flag~2_combout ),
	.datae(!\aempty_flag~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~4 .extended_lut = "off";
defparam \aempty_flag~4 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \aempty_flag~4 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~5 (
	.dataa(!\LessThan3~0_combout ),
	.datab(!\LessThan3~7_combout ),
	.datac(!\LessThan3~8_combout ),
	.datad(!\aempty_flag~0_combout ),
	.datae(!\aempty_flag~1_combout ),
	.dataf(!\aempty_flag~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~5 .extended_lut = "off";
defparam \aempty_flag~5 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \aempty_flag~5 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_5 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_0,
	g_out_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	g_out_10;
input 	g_out_9;
input 	g_out_8;
input 	g_out_7;
input 	g_out_6;
input 	g_out_5;
input 	g_out_4;
input 	g_out_3;
input 	g_out_2;
input 	g_out_0;
input 	g_out_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_78 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.g_out_7(g_out_7),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_77 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.g_out_6(g_out_6),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_76 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.g_out_5(g_out_5),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_75 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.g_out_4(g_out_4),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_74 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.g_out_3(g_out_3),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_71 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.g_out_10(g_out_10),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_80 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.g_out_9(g_out_9),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_79 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.g_out_8(g_out_8),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_73 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.g_out_2(g_out_2),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_72 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.g_out_1(g_out_1),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_70 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.g_out_0(g_out_0),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_70 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_0,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_0;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_70 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_0),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_70 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_71 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_10,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_10;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_71 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_10),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_71 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_72 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_72 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_72 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_73 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_2,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_2;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_73 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_2),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_73 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_74 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_3,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_3;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_74 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_3),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_74 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_75 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_4,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_4;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_75 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_4),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_75 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_76 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_5,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_5;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_76 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_5),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_76 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_77 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_6,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_6;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_77 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_6),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_77 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_78 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_7,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_7;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_78 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_7),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_78 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_79 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_8,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_8;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_79 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_8),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_79 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_80 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_9,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_9;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_80 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_9),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_80 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_6 (
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_82 \sync[10].u (
	.dreg_1(dreg_1),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_91 \sync[9].u (
	.dreg_1(dreg_19),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_90 \sync[8].u (
	.dreg_1(dreg_110),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_89 \sync[7].u (
	.dreg_1(dreg_17),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_88 \sync[6].u (
	.dreg_1(dreg_18),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_87 \sync[5].u (
	.dreg_1(dreg_15),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_86 \sync[4].u (
	.dreg_1(dreg_16),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_85 \sync[3].u (
	.dreg_1(dreg_13),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_84 \sync[2].u (
	.dreg_1(dreg_14),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_83 \sync[1].u (
	.dreg_1(dreg_12),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_81 \sync[0].u (
	.dreg_1(dreg_11),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_81 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_81 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_81 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_82 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_82 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_82 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_83 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_83 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_83 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_84 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_84 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_84 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_85 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_85 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_85 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_86 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_86 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_86 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_87 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_87 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_87 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_88 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_88 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_88 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_89 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_89 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_89 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_90 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_90 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_90 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_91 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_91 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_91 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_7 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	g_out_10;
input 	g_out_9;
input 	g_out_8;
input 	g_out_7;
input 	g_out_6;
input 	g_out_5;
input 	g_out_4;
input 	g_out_3;
input 	g_out_2;
input 	g_out_1;
input 	g_out_0;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_93 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.g_out_10(g_out_10),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_102 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.g_out_9(g_out_9),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_101 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.g_out_8(g_out_8),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_100 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.g_out_7(g_out_7),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_99 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.g_out_6(g_out_6),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_98 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.g_out_5(g_out_5),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_97 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.g_out_4(g_out_4),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_96 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.g_out_3(g_out_3),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_95 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.g_out_2(g_out_2),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_94 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.g_out_1(g_out_1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_92 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.g_out_0(g_out_0),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_92 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_0,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_0;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_92 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_0),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_92 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_93 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_10,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_10;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_93 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_10),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_93 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_94 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_94 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_94 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_95 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_2,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_2;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_95 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_2),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_95 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_96 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_3,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_3;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_96 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_3),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_96 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_97 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_4,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_4;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_97 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_4),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_97 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_98 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_5,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_5;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_98 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_5),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_98 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_99 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_6,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_6;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_99 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_6),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_99 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_100 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_7,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_7;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_100 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_7),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_100 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_101 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_8,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_8;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_101 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_8),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_101 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_102 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_9,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_9;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_102 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_9),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_102 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_8 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_104 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_113 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_108 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_107 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_106 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_105 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_103 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_112 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_111 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_110 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_109 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_103 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_103 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_103 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_104 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_104 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_104 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_105 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_105 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_105 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_106 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_106 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_106 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_107 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_107 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_107 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_108 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_108 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_108 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_109 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_109 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_109 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_110 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_110 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_110 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_111 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_111 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_111 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_112 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_112 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_112 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_113 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_113 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_113 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_1 (
	q_b_32,
	q_b_39,
	q_b_34,
	q_b_33,
	q_b_36,
	q_b_35,
	q_b_37,
	rx_wren32,
	rx_eop32,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	b_out_9,
	b_out_10,
	b_out_01,
	b_out_11,
	b_out_21,
	b_out_31,
	b_out_41,
	b_out_51,
	b_out_61,
	b_out_71,
	b_out_81,
	b_out_91,
	b_out_101,
	byte_empty_1,
	frm_type32_0,
	rx_sop32,
	frm_type32_2,
	frm_type32_1,
	GND_port,
	clk_32_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_32;
output 	q_b_39;
output 	q_b_34;
output 	q_b_33;
output 	q_b_36;
output 	q_b_35;
output 	q_b_37;
input 	rx_wren32;
input 	rx_eop32;
input 	b_out_0;
input 	b_out_1;
input 	b_out_2;
input 	b_out_3;
input 	b_out_4;
input 	b_out_5;
input 	b_out_6;
input 	b_out_7;
input 	b_out_8;
input 	b_out_9;
input 	b_out_10;
input 	b_out_01;
input 	b_out_11;
input 	b_out_21;
input 	b_out_31;
input 	b_out_41;
input 	b_out_51;
input 	b_out_61;
input 	b_out_71;
input 	b_out_81;
input 	b_out_91;
input 	b_out_101;
input 	byte_empty_1;
input 	frm_type32_0;
input 	rx_sop32;
input 	frm_type32_2;
input 	frm_type32_1;
input 	GND_port;
input 	clk_32_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_3 altsyncram_component(
	.q_b({q_b_39,q_b_unconnected_wire_38,q_b_37,q_b_36,q_b_35,q_b_34,q_b_33,q_b_32,q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,
q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,
q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,
q_b_unconnected_wire_1,q_b_unconnected_wire_0}),
	.wren_a(rx_wren32),
	.data_a({byte_empty_1,gnd,GND_port,frm_type32_2,frm_type32_1,frm_type32_0,rx_sop32,rx_eop32,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.address_a({b_out_10,b_out_9,b_out_8,b_out_7,b_out_6,b_out_5,b_out_4,b_out_3,b_out_2,b_out_1,b_out_0}),
	.address_b({b_out_101,b_out_91,b_out_81,b_out_71,b_out_61,b_out_51,b_out_41,b_out_31,b_out_21,b_out_11,b_out_01}),
	.clock1(clk_32_clk),
	.clock0(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altsyncram_3 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	wren_a;
input 	[39:0] data_a;
input 	[10:0] address_a;
input 	[10:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_p9o1 auto_generated(
	.q_b({q_b[39],q_b_unconnected_wire_38,q_b[37],q_b[36],q_b[35],q_b[34],q_b[33],q_b[32],q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,
q_b_unconnected_wire_22,q_b_unconnected_wire_21,q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,
q_b_unconnected_wire_11,q_b_unconnected_wire_10,q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_unconnected_wire_1,
q_b_unconnected_wire_0}),
	.wren_a(wren_a),
	.data_a({data_a[39],gnd,data_a[37],data_a[36],data_a[35],data_a[34],data_a[33],data_a[32],gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.address_a({address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock1(clock1),
	.clock0(clock0));

endmodule

module IoTOctopus_QSYS_altsyncram_p9o1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	wren_a;
input 	[39:0] data_a;
input 	[10:0] address_a;
input 	[10:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a39_PORTBDATAOUT_bus;
wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;

assign q_b[32] = ram_block1a32_PORTBDATAOUT_bus[0];

assign q_b[39] = ram_block1a39_PORTBDATAOUT_bus[0];

assign q_b[34] = ram_block1a34_PORTBDATAOUT_bus[0];

assign q_b[33] = ram_block1a33_PORTBDATAOUT_bus[0];

assign q_b[36] = ram_block1a36_PORTBDATAOUT_bus[0];

assign q_b[35] = ram_block1a35_PORTBDATAOUT_bus[0];

assign q_b[37] = ram_block1a37_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a32(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 11;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 2047;
defparam ram_block1a32.port_a_logical_ram_depth = 2048;
defparam ram_block1a32.port_a_logical_ram_width = 40;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 11;
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "none";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 2047;
defparam ram_block1a32.port_b_logical_ram_depth = 2048;
defparam ram_block1a32.port_b_logical_ram_width = 40;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";

cyclonev_ram_block ram_block1a39(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[39]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a39_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a39.operation_mode = "dual_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 11;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 0;
defparam ram_block1a39.port_a_first_bit_number = 39;
defparam ram_block1a39.port_a_last_address = 2047;
defparam ram_block1a39.port_a_logical_ram_depth = 2048;
defparam ram_block1a39.port_a_logical_ram_width = 40;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_address_clear = "none";
defparam ram_block1a39.port_b_address_clock = "clock1";
defparam ram_block1a39.port_b_address_width = 11;
defparam ram_block1a39.port_b_data_out_clear = "none";
defparam ram_block1a39.port_b_data_out_clock = "none";
defparam ram_block1a39.port_b_data_width = 1;
defparam ram_block1a39.port_b_first_address = 0;
defparam ram_block1a39.port_b_first_bit_number = 39;
defparam ram_block1a39.port_b_last_address = 2047;
defparam ram_block1a39.port_b_logical_ram_depth = 2048;
defparam ram_block1a39.port_b_logical_ram_width = 40;
defparam ram_block1a39.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a39.port_b_read_enable_clock = "clock1";
defparam ram_block1a39.ram_block_type = "auto";

cyclonev_ram_block ram_block1a34(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 11;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 2047;
defparam ram_block1a34.port_a_logical_ram_depth = 2048;
defparam ram_block1a34.port_a_logical_ram_width = 40;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 11;
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "none";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 2047;
defparam ram_block1a34.port_b_logical_ram_depth = 2048;
defparam ram_block1a34.port_b_logical_ram_width = 40;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";

cyclonev_ram_block ram_block1a33(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 11;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 2047;
defparam ram_block1a33.port_a_logical_ram_depth = 2048;
defparam ram_block1a33.port_a_logical_ram_width = 40;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 11;
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "none";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 2047;
defparam ram_block1a33.port_b_logical_ram_depth = 2048;
defparam ram_block1a33.port_b_logical_ram_width = 40;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";

cyclonev_ram_block ram_block1a36(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 11;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 0;
defparam ram_block1a36.port_a_first_bit_number = 36;
defparam ram_block1a36.port_a_last_address = 2047;
defparam ram_block1a36.port_a_logical_ram_depth = 2048;
defparam ram_block1a36.port_a_logical_ram_width = 40;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 11;
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "none";
defparam ram_block1a36.port_b_data_width = 1;
defparam ram_block1a36.port_b_first_address = 0;
defparam ram_block1a36.port_b_first_bit_number = 36;
defparam ram_block1a36.port_b_last_address = 2047;
defparam ram_block1a36.port_b_logical_ram_depth = 2048;
defparam ram_block1a36.port_b_logical_ram_width = 40;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";

cyclonev_ram_block ram_block1a35(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 11;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 2047;
defparam ram_block1a35.port_a_logical_ram_depth = 2048;
defparam ram_block1a35.port_a_logical_ram_width = 40;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 11;
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "none";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 2047;
defparam ram_block1a35.port_b_logical_ram_depth = 2048;
defparam ram_block1a35.port_b_logical_ram_width = 40;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";

cyclonev_ram_block ram_block1a37(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_rx_min_ff:U_RXFF|altera_tse_a_fifo_opt_1246:RX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_p9o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 11;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 0;
defparam ram_block1a37.port_a_first_bit_number = 37;
defparam ram_block1a37.port_a_last_address = 2047;
defparam ram_block1a37.port_a_logical_ram_depth = 2048;
defparam ram_block1a37.port_a_logical_ram_width = 40;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 11;
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "none";
defparam ram_block1a37.port_b_data_width = 1;
defparam ram_block1a37.port_b_first_address = 0;
defparam ram_block1a37.port_b_first_bit_number = 37;
defparam ram_block1a37.port_b_last_address = 2047;
defparam ram_block1a37.port_b_logical_ram_depth = 2048;
defparam ram_block1a37.port_b_logical_ram_width = 40;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_3 (
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	b_out_9,
	b_out_10,
	reset,
	data_rdreq,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_0,
	g_out_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	b_out_5;
output 	b_out_6;
output 	b_out_7;
output 	b_out_8;
output 	b_out_9;
output 	b_out_10;
input 	reset;
input 	data_rdreq;
output 	g_out_10;
output 	g_out_9;
output 	g_out_8;
output 	g_out_7;
output 	g_out_6;
output 	g_out_5;
output 	g_out_4;
output 	g_out_3;
output 	g_out_2;
output 	g_out_0;
output 	g_out_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \b_int[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \b_int[3]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \b_int[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \b_int[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \b_int[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \b_int[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \b_int[8]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \b_int[9]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \b_int[10]~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \b_int[1]~q ;
wire \Add0~1_sumout ;
wire \b_int~0_combout ;
wire \b_int[0]~q ;
wire \b_out[0]~0_combout ;
wire \gry_grayval[9]~combout ;
wire \gry_grayval[8]~combout ;
wire \gry_grayval[7]~combout ;
wire \gry_grayval[6]~combout ;
wire \gry_grayval[5]~combout ;
wire \gry_grayval[4]~combout ;
wire \gry_grayval[3]~combout ;
wire \gry_grayval[2]~combout ;
wire \gry_grayval[0]~combout ;
wire \gry_grayval[1]~combout ;


dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[5] (
	.clk(clk),
	.d(\b_int[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[6] (
	.clk(clk),
	.d(\b_int[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[7] (
	.clk(clk),
	.d(\b_int[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

dffeas \b_out[9] (
	.clk(clk),
	.d(\b_int[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_9),
	.prn(vcc));
defparam \b_out[9] .is_wysiwyg = "true";
defparam \b_out[9] .power_up = "low";

dffeas \b_out[10] (
	.clk(clk),
	.d(\b_int[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(b_out_10),
	.prn(vcc));
defparam \b_out[10] .is_wysiwyg = "true";
defparam \b_out[10] .power_up = "low";

dffeas \g_out[10] (
	.clk(clk),
	.d(\b_int[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_10),
	.prn(vcc));
defparam \g_out[10] .is_wysiwyg = "true";
defparam \g_out[10] .power_up = "low";

dffeas \g_out[9] (
	.clk(clk),
	.d(\gry_grayval[9]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_9),
	.prn(vcc));
defparam \g_out[9] .is_wysiwyg = "true";
defparam \g_out[9] .power_up = "low";

dffeas \g_out[8] (
	.clk(clk),
	.d(\gry_grayval[8]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_8),
	.prn(vcc));
defparam \g_out[8] .is_wysiwyg = "true";
defparam \g_out[8] .power_up = "low";

dffeas \g_out[7] (
	.clk(clk),
	.d(\gry_grayval[7]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_7),
	.prn(vcc));
defparam \g_out[7] .is_wysiwyg = "true";
defparam \g_out[7] .power_up = "low";

dffeas \g_out[6] (
	.clk(clk),
	.d(\gry_grayval[6]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_6),
	.prn(vcc));
defparam \g_out[6] .is_wysiwyg = "true";
defparam \g_out[6] .power_up = "low";

dffeas \g_out[5] (
	.clk(clk),
	.d(\gry_grayval[5]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_5),
	.prn(vcc));
defparam \g_out[5] .is_wysiwyg = "true";
defparam \g_out[5] .power_up = "low";

dffeas \g_out[4] (
	.clk(clk),
	.d(\gry_grayval[4]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[3] (
	.clk(clk),
	.d(\gry_grayval[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[2] (
	.clk(clk),
	.d(\gry_grayval[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[0] (
	.clk(clk),
	.d(\gry_grayval[0]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

dffeas \g_out[1] (
	.clk(clk),
	.d(\gry_grayval[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \b_int[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \b_int[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[5]~q ),
	.prn(vcc));
defparam \b_int[5] .is_wysiwyg = "true";
defparam \b_int[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \b_int[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[6]~q ),
	.prn(vcc));
defparam \b_int[6] .is_wysiwyg = "true";
defparam \b_int[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \b_int[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[7]~q ),
	.prn(vcc));
defparam \b_int[7] .is_wysiwyg = "true";
defparam \b_int[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \b_int[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[8]~q ),
	.prn(vcc));
defparam \b_int[8] .is_wysiwyg = "true";
defparam \b_int[8] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \b_int[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[9]~q ),
	.prn(vcc));
defparam \b_int[9] .is_wysiwyg = "true";
defparam \b_int[9] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \b_int[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[10]~q ),
	.prn(vcc));
defparam \b_int[10] .is_wysiwyg = "true";
defparam \b_int[10] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[5]~q ),
	.datac(!\b_int[8]~q ),
	.datad(!\b_int[9]~q ),
	.datae(!\b_int[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[3]~q ),
	.datac(!\b_int[4]~q ),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[7]~q ),
	.datac(!\LessThan0~0_combout ),
	.datad(!\LessThan0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~2 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \b_int~0 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[7]~q ),
	.datac(!\Add0~1_sumout ),
	.datad(!\LessThan0~0_combout ),
	.datae(!\LessThan0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int~0 .extended_lut = "off";
defparam \b_int~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \b_int~0 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(data_rdreq),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[9] (
	.dataa(!\b_int[9]~q ),
	.datab(!\b_int[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[9] .extended_lut = "off";
defparam \gry_grayval[9] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[9] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[8] (
	.dataa(!\b_int[8]~q ),
	.datab(!\b_int[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[8] .extended_lut = "off";
defparam \gry_grayval[8] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[8] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[7] (
	.dataa(!\b_int[7]~q ),
	.datab(!\b_int[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[7] .extended_lut = "off";
defparam \gry_grayval[7] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[7] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[6] (
	.dataa(!\b_int[6]~q ),
	.datab(!\b_int[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[6] .extended_lut = "off";
defparam \gry_grayval[6] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[6] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[5] (
	.dataa(!\b_int[5]~q ),
	.datab(!\b_int[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[5] .extended_lut = "off";
defparam \gry_grayval[5] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[5] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[4] (
	.dataa(!\b_int[4]~q ),
	.datab(!\b_int[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[4] .extended_lut = "off";
defparam \gry_grayval[4] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[4] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[3] (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[3] .extended_lut = "off";
defparam \gry_grayval[3] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[3] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[2] (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[2] .extended_lut = "off";
defparam \gry_grayval[2] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[2] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[0] (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[0] .extended_lut = "off";
defparam \gry_grayval[0] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[0] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[1] (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[1] .extended_lut = "off";
defparam \gry_grayval[1] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[1] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_4 (
	rx_wren32,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	b_out_9,
	b_out_10,
	reset,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rx_wren32;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	b_out_5;
output 	b_out_6;
output 	b_out_7;
output 	b_out_8;
output 	b_out_9;
output 	b_out_10;
input 	reset;
output 	g_out_10;
output 	g_out_9;
output 	g_out_8;
output 	g_out_7;
output 	g_out_6;
output 	g_out_5;
output 	g_out_4;
output 	g_out_3;
output 	g_out_2;
output 	g_out_1;
output 	g_out_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \b_int[2]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \b_int[3]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \b_int[4]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \b_int[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \b_int[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \b_int[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \b_int[8]~q ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \b_int[9]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \b_int[10]~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \b_int[1]~q ;
wire \Add0~1_sumout ;
wire \b_int~0_combout ;
wire \b_int[0]~q ;
wire \b_out[0]~0_combout ;
wire \gry_grayval[9]~combout ;
wire \gry_grayval[8]~combout ;
wire \gry_grayval[7]~combout ;
wire \gry_grayval[6]~combout ;
wire \gry_grayval[5]~combout ;
wire \gry_grayval[4]~combout ;
wire \gry_grayval[3]~combout ;
wire \gry_grayval[2]~combout ;
wire \gry_grayval[1]~combout ;
wire \gry_grayval[0]~combout ;


dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[5] (
	.clk(clk),
	.d(\b_int[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[6] (
	.clk(clk),
	.d(\b_int[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[7] (
	.clk(clk),
	.d(\b_int[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

dffeas \b_out[9] (
	.clk(clk),
	.d(\b_int[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_9),
	.prn(vcc));
defparam \b_out[9] .is_wysiwyg = "true";
defparam \b_out[9] .power_up = "low";

dffeas \b_out[10] (
	.clk(clk),
	.d(\b_int[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(b_out_10),
	.prn(vcc));
defparam \b_out[10] .is_wysiwyg = "true";
defparam \b_out[10] .power_up = "low";

dffeas \g_out[10] (
	.clk(clk),
	.d(\b_int[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_10),
	.prn(vcc));
defparam \g_out[10] .is_wysiwyg = "true";
defparam \g_out[10] .power_up = "low";

dffeas \g_out[9] (
	.clk(clk),
	.d(\gry_grayval[9]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_9),
	.prn(vcc));
defparam \g_out[9] .is_wysiwyg = "true";
defparam \g_out[9] .power_up = "low";

dffeas \g_out[8] (
	.clk(clk),
	.d(\gry_grayval[8]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_8),
	.prn(vcc));
defparam \g_out[8] .is_wysiwyg = "true";
defparam \g_out[8] .power_up = "low";

dffeas \g_out[7] (
	.clk(clk),
	.d(\gry_grayval[7]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_7),
	.prn(vcc));
defparam \g_out[7] .is_wysiwyg = "true";
defparam \g_out[7] .power_up = "low";

dffeas \g_out[6] (
	.clk(clk),
	.d(\gry_grayval[6]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_6),
	.prn(vcc));
defparam \g_out[6] .is_wysiwyg = "true";
defparam \g_out[6] .power_up = "low";

dffeas \g_out[5] (
	.clk(clk),
	.d(\gry_grayval[5]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_5),
	.prn(vcc));
defparam \g_out[5] .is_wysiwyg = "true";
defparam \g_out[5] .power_up = "low";

dffeas \g_out[4] (
	.clk(clk),
	.d(\gry_grayval[4]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[3] (
	.clk(clk),
	.d(\gry_grayval[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[2] (
	.clk(clk),
	.d(\gry_grayval[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[1] (
	.clk(clk),
	.d(\gry_grayval[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[0] (
	.clk(clk),
	.d(\gry_grayval[0]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \b_int[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \b_int[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[5]~q ),
	.prn(vcc));
defparam \b_int[5] .is_wysiwyg = "true";
defparam \b_int[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \b_int[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[6]~q ),
	.prn(vcc));
defparam \b_int[6] .is_wysiwyg = "true";
defparam \b_int[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \b_int[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[7]~q ),
	.prn(vcc));
defparam \b_int[7] .is_wysiwyg = "true";
defparam \b_int[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \b_int[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[8]~q ),
	.prn(vcc));
defparam \b_int[8] .is_wysiwyg = "true";
defparam \b_int[8] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \b_int[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[9]~q ),
	.prn(vcc));
defparam \b_int[9] .is_wysiwyg = "true";
defparam \b_int[9] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \b_int[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[10]~q ),
	.prn(vcc));
defparam \b_int[10] .is_wysiwyg = "true";
defparam \b_int[10] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[2]~q ),
	.datac(!\b_int[8]~q ),
	.datad(!\b_int[9]~q ),
	.datae(!\b_int[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(!\b_int[5]~q ),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[7]~q ),
	.datac(!\LessThan0~0_combout ),
	.datad(!\LessThan0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~2 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \b_int~0 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[7]~q ),
	.datac(!\Add0~1_sumout ),
	.datad(!\LessThan0~0_combout ),
	.datae(!\LessThan0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int~0 .extended_lut = "off";
defparam \b_int~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \b_int~0 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rx_wren32),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[9] (
	.dataa(!\b_int[9]~q ),
	.datab(!\b_int[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[9] .extended_lut = "off";
defparam \gry_grayval[9] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[9] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[8] (
	.dataa(!\b_int[8]~q ),
	.datab(!\b_int[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[8] .extended_lut = "off";
defparam \gry_grayval[8] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[8] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[7] (
	.dataa(!\b_int[7]~q ),
	.datab(!\b_int[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[7] .extended_lut = "off";
defparam \gry_grayval[7] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[7] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[6] (
	.dataa(!\b_int[6]~q ),
	.datab(!\b_int[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[6] .extended_lut = "off";
defparam \gry_grayval[6] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[6] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[5] (
	.dataa(!\b_int[5]~q ),
	.datab(!\b_int[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[5] .extended_lut = "off";
defparam \gry_grayval[5] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[5] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[4] (
	.dataa(!\b_int[4]~q ),
	.datab(!\b_int[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[4] .extended_lut = "off";
defparam \gry_grayval[4] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[4] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[3] (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[3] .extended_lut = "off";
defparam \gry_grayval[3] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[3] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[2] (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[2] .extended_lut = "off";
defparam \gry_grayval[2] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[2] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[1] (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[1] .extended_lut = "off";
defparam \gry_grayval[1] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[1] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[0] (
	.dataa(!\b_int[0]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[0] .extended_lut = "off";
defparam \gry_grayval[0] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[0] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_top_1geth (
	q_b_9,
	eop_sft_0,
	q_b_8,
	en,
	data_3,
	data_2,
	data_1,
	data_0,
	data_7,
	data_6,
	data_5,
	data_4,
	q_b_4,
	dout_reg_sft_28,
	q_b_0,
	dout_reg_sft_24,
	q_b_5,
	dout_reg_sft_29,
	q_b_1,
	dout_reg_sft_25,
	q_b_6,
	dout_reg_sft_30,
	q_b_2,
	dout_reg_sft_26,
	q_b_7,
	dout_reg_sft_31,
	q_b_3,
	dout_reg_sft_27,
	err,
	tx_ff_uflow,
	afull_flag,
	txclk_ena,
	altera_tse_reset_synchronizer_chain_out,
	rx_stat_wren,
	payload_length_0,
	payload_length_1,
	payload_length_2,
	payload_length_3,
	payload_length_4,
	payload_length_5,
	payload_length_6,
	payload_length_7,
	payload_length_8,
	payload_length_9,
	payload_length_10,
	payload_length_11,
	payload_length_12,
	payload_length_13,
	payload_length_14,
	payload_length_15,
	altera_tse_reset_synchronizer_chain_out1,
	tx_empty,
	tx_data_int_7,
	dreg_1,
	tx_en_s_1,
	rxclk_ena,
	rx_wren_int,
	rx_eop_int,
	rx_stat_data_s_5,
	rx_stat_data_s_0,
	rx_stat_data_s_1,
	rx_stat_data_s_2,
	rx_stat_data_s_3,
	rx_sop_int,
	rx_ucast,
	rx_mcast,
	rx_bcast,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err,
	tx_eop_int,
	empty_flag,
	always9,
	col_int,
	always91,
	tx_rden_mii,
	tx_rden_int,
	always92,
	mac_ena,
	sav_flag,
	rx_data_val,
	magic_pkt_ena,
	ethernet_mode,
	dreg_11,
	tx_stat_1,
	rx_done_reg,
	sop_reg,
	tx_stat_rden,
	sleep_ena,
	rx_data_int_3,
	rx_data_int_2,
	rx_data_int_1,
	rx_data_int_0,
	rx_data_int_7,
	rx_data_int_6,
	rx_data_int_5,
	rx_data_int_4,
	dreg_12,
	m_rx_crs,
	tx_stat_0,
	GND_port,
	mac_tx_clock_connection_clk,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	q_b_9;
input 	eop_sft_0;
input 	q_b_8;
input 	en;
input 	data_3;
input 	data_2;
input 	data_1;
input 	data_0;
input 	data_7;
input 	data_6;
input 	data_5;
input 	data_4;
input 	q_b_4;
input 	dout_reg_sft_28;
input 	q_b_0;
input 	dout_reg_sft_24;
input 	q_b_5;
input 	dout_reg_sft_29;
input 	q_b_1;
input 	dout_reg_sft_25;
input 	q_b_6;
input 	dout_reg_sft_30;
input 	q_b_2;
input 	dout_reg_sft_26;
input 	q_b_7;
input 	dout_reg_sft_31;
input 	q_b_3;
input 	dout_reg_sft_27;
input 	err;
output 	tx_ff_uflow;
input 	afull_flag;
input 	txclk_ena;
input 	altera_tse_reset_synchronizer_chain_out;
output 	rx_stat_wren;
output 	payload_length_0;
output 	payload_length_1;
output 	payload_length_2;
output 	payload_length_3;
output 	payload_length_4;
output 	payload_length_5;
output 	payload_length_6;
output 	payload_length_7;
output 	payload_length_8;
output 	payload_length_9;
output 	payload_length_10;
output 	payload_length_11;
output 	payload_length_12;
output 	payload_length_13;
output 	payload_length_14;
output 	payload_length_15;
input 	altera_tse_reset_synchronizer_chain_out1;
input 	tx_empty;
input 	tx_data_int_7;
output 	dreg_1;
output 	tx_en_s_1;
input 	rxclk_ena;
output 	rx_wren_int;
output 	rx_eop_int;
output 	rx_stat_data_s_5;
output 	rx_stat_data_s_0;
output 	rx_stat_data_s_1;
output 	rx_stat_data_s_2;
output 	rx_stat_data_s_3;
output 	rx_sop_int;
output 	rx_ucast;
output 	rx_mcast;
output 	rx_bcast;
output 	rd_14_4;
output 	rd_14_0;
output 	rd_14_5;
output 	rd_14_1;
output 	rd_14_6;
output 	rd_14_2;
output 	rd_14_7;
output 	rd_14_3;
output 	tx_err;
input 	tx_eop_int;
input 	empty_flag;
output 	always9;
output 	col_int;
output 	always91;
output 	tx_rden_mii;
output 	tx_rden_int;
output 	always92;
input 	mac_ena;
input 	sav_flag;
output 	rx_data_val;
output 	magic_pkt_ena;
input 	ethernet_mode;
output 	dreg_11;
input 	tx_stat_1;
output 	rx_done_reg;
input 	sop_reg;
output 	tx_stat_rden;
input 	sleep_ena;
output 	rx_data_int_3;
output 	rx_data_int_2;
output 	rx_data_int_1;
output 	rx_data_int_0;
output 	rx_data_int_7;
output 	rx_data_int_6;
output 	rx_data_int_5;
output 	rx_data_int_4;
input 	dreg_12;
input 	m_rx_crs;
input 	tx_stat_0;
input 	GND_port;
input 	mac_tx_clock_connection_clk;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_tse_mac_tx U_TX(
	.q_b_9(q_b_9),
	.eop_sft_0(eop_sft_0),
	.q_b_8(q_b_8),
	.q_b_4(q_b_4),
	.dout_reg_sft_28(dout_reg_sft_28),
	.q_b_0(q_b_0),
	.dout_reg_sft_24(dout_reg_sft_24),
	.q_b_5(q_b_5),
	.dout_reg_sft_29(dout_reg_sft_29),
	.q_b_1(q_b_1),
	.dout_reg_sft_25(dout_reg_sft_25),
	.q_b_6(q_b_6),
	.dout_reg_sft_30(dout_reg_sft_30),
	.q_b_2(q_b_2),
	.dout_reg_sft_26(dout_reg_sft_26),
	.q_b_7(q_b_7),
	.dout_reg_sft_31(dout_reg_sft_31),
	.q_b_3(q_b_3),
	.dout_reg_sft_27(dout_reg_sft_27),
	.tx_ff_uflow1(tx_ff_uflow),
	.txclk_ena(txclk_ena),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.tx_empty(tx_empty),
	.tx_data_int_7(tx_data_int_7),
	.dreg_1(dreg_1),
	.tx_en_s_1(tx_en_s_1),
	.rd_14_4(rd_14_4),
	.rd_14_0(rd_14_0),
	.rd_14_5(rd_14_5),
	.rd_14_1(rd_14_1),
	.rd_14_6(rd_14_6),
	.rd_14_2(rd_14_2),
	.rd_14_7(rd_14_7),
	.rd_14_3(rd_14_3),
	.tx_err1(tx_err),
	.tx_eop_int(tx_eop_int),
	.empty_flag(empty_flag),
	.always9(always9),
	.col_int1(col_int),
	.always91(always91),
	.tx_rden_mii1(tx_rden_mii),
	.tx_rden_int(tx_rden_int),
	.always92(always92),
	.mac_ena(mac_ena),
	.tx_sav_int(sav_flag),
	.ethernet_mode(ethernet_mode),
	.dreg_11(dreg_11),
	.tx_stat_1(tx_stat_1),
	.sop_reg(sop_reg),
	.tx_stat_rden1(tx_stat_rden),
	.sleep_ena(sleep_ena),
	.dreg_12(dreg_12),
	.m_rx_crs(m_rx_crs),
	.tx_stat_0(tx_stat_0),
	.GND_port(GND_port),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_mac_rx U_RX(
	.en(en),
	.rx_d({data_7,data_6,data_5,data_4,data_3,data_2,data_1,data_0}),
	.err(err),
	.afull_flag(afull_flag),
	.rx_stat_wren1(rx_stat_wren),
	.payload_length_0(payload_length_0),
	.payload_length_1(payload_length_1),
	.payload_length_2(payload_length_2),
	.payload_length_3(payload_length_3),
	.payload_length_4(payload_length_4),
	.payload_length_5(payload_length_5),
	.payload_length_6(payload_length_6),
	.payload_length_7(payload_length_7),
	.payload_length_8(payload_length_8),
	.payload_length_9(payload_length_9),
	.payload_length_10(payload_length_10),
	.payload_length_11(payload_length_11),
	.payload_length_12(payload_length_12),
	.payload_length_13(payload_length_13),
	.payload_length_14(payload_length_14),
	.payload_length_15(payload_length_15),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.rxclk_ena(rxclk_ena),
	.rx_wren_int1(rx_wren_int),
	.rx_eop_int1(rx_eop_int),
	.rx_stat_data_s_5(rx_stat_data_s_5),
	.rx_stat_data_s_0(rx_stat_data_s_0),
	.rx_stat_data_s_1(rx_stat_data_s_1),
	.rx_stat_data_s_2(rx_stat_data_s_2),
	.rx_stat_data_s_3(rx_stat_data_s_3),
	.rx_sop_int1(rx_sop_int),
	.rx_ucast1(rx_ucast),
	.rx_mcast1(rx_mcast),
	.rx_bcast1(rx_bcast),
	.rx_data_val1(rx_data_val),
	.magic_pkt_ena1(magic_pkt_ena),
	.ethernet_mode(ethernet_mode),
	.rx_done_reg1(rx_done_reg),
	.sleep_ena(sleep_ena),
	.rx_data_int_3(rx_data_int_3),
	.rx_data_int_2(rx_data_int_2),
	.rx_data_int_1(rx_data_int_1),
	.rx_data_int_0(rx_data_int_0),
	.rx_data_int_7(rx_data_int_7),
	.rx_data_int_6(rx_data_int_6),
	.rx_data_int_5(rx_data_int_5),
	.rx_data_int_4(rx_data_int_4),
	.dreg_1(dreg_12),
	.GND_port(GND_port),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_tse_mac_rx (
	en,
	rx_d,
	err,
	afull_flag,
	rx_stat_wren1,
	payload_length_0,
	payload_length_1,
	payload_length_2,
	payload_length_3,
	payload_length_4,
	payload_length_5,
	payload_length_6,
	payload_length_7,
	payload_length_8,
	payload_length_9,
	payload_length_10,
	payload_length_11,
	payload_length_12,
	payload_length_13,
	payload_length_14,
	payload_length_15,
	altera_tse_reset_synchronizer_chain_out,
	rxclk_ena,
	rx_wren_int1,
	rx_eop_int1,
	rx_stat_data_s_5,
	rx_stat_data_s_0,
	rx_stat_data_s_1,
	rx_stat_data_s_2,
	rx_stat_data_s_3,
	rx_sop_int1,
	rx_ucast1,
	rx_mcast1,
	rx_bcast1,
	rx_data_val1,
	magic_pkt_ena1,
	ethernet_mode,
	rx_done_reg1,
	sleep_ena,
	rx_data_int_3,
	rx_data_int_2,
	rx_data_int_1,
	rx_data_int_0,
	rx_data_int_7,
	rx_data_int_6,
	rx_data_int_5,
	rx_data_int_4,
	dreg_1,
	GND_port,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	en;
input 	[7:0] rx_d;
input 	err;
input 	afull_flag;
output 	rx_stat_wren1;
output 	payload_length_0;
output 	payload_length_1;
output 	payload_length_2;
output 	payload_length_3;
output 	payload_length_4;
output 	payload_length_5;
output 	payload_length_6;
output 	payload_length_7;
output 	payload_length_8;
output 	payload_length_9;
output 	payload_length_10;
output 	payload_length_11;
output 	payload_length_12;
output 	payload_length_13;
output 	payload_length_14;
output 	payload_length_15;
input 	altera_tse_reset_synchronizer_chain_out;
input 	rxclk_ena;
output 	rx_wren_int1;
output 	rx_eop_int1;
output 	rx_stat_data_s_5;
output 	rx_stat_data_s_0;
output 	rx_stat_data_s_1;
output 	rx_stat_data_s_2;
output 	rx_stat_data_s_3;
output 	rx_sop_int1;
output 	rx_ucast1;
output 	rx_mcast1;
output 	rx_bcast1;
output 	rx_data_val1;
output 	magic_pkt_ena1;
input 	ethernet_mode;
output 	rx_done_reg1;
input 	sleep_ena;
output 	rx_data_int_3;
output 	rx_data_int_2;
output 	rx_data_int_1;
output 	rx_data_int_0;
output 	rx_data_int_7;
output 	rx_data_int_6;
output 	rx_data_int_5;
output 	rx_data_int_4;
input 	dreg_1;
input 	GND_port;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout ;
wire \U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ;
wire \U_SYNC_2|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_11|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_7|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_6|std_sync_no_cut|dreg[1]~q ;
wire \U_CRC|eof_dly[2]~q ;
wire \U_CRC|crc_ok~q ;
wire \U_SYNC_4|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_PAD_ENA|std_sync_no_cut|dreg[1]~q ;
wire \eof_crc~0_combout ;
wire \U_SYNC_9|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_10|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_13|std_sync_no_cut|dreg[1]~q ;
wire \enable_rx_reg3~0_combout ;
wire \enable_rx_reg3~q ;
wire \rx_en_s~0_combout ;
wire \rx_en_s[0]~q ;
wire \rx_en_s[1]~q ;
wire \rx_en_s[2]~q ;
wire \rx_en_s[3]~q ;
wire \rx_en_s[4]~q ;
wire \rx_en_s[5]~q ;
wire \rx_en_s[6]~q ;
wire \rx_en_s[7]~q ;
wire \rx_en_s[8]~q ;
wire \rx_en_s[9]~q ;
wire \rx_en_s[10]~q ;
wire \rx_en_s[11]~q ;
wire \rx_en_s[12]~q ;
wire \rx_en_s[13]~q ;
wire \rx_en_s[14]~q ;
wire \rx_en_s[15]~q ;
wire \rx_en_s[16]~q ;
wire \rx_en_s[17]~q ;
wire \rx_en_s[18]~q ;
wire \rx_en_s[19]~q ;
wire \rx_en_s[20]~q ;
wire \rx_en_s[21]~q ;
wire \rx_en_s[22]~q ;
wire \rx_en_s[23]~q ;
wire \rx_en_s[24]~q ;
wire \rxd_0[0]~q ;
wire \rxd_1[0]~q ;
wire \rxd_2[0]~q ;
wire \rxd_3[0]~q ;
wire \rxd_4[0]~q ;
wire \rxd_5[0]~q ;
wire \rxd_6[0]~q ;
wire \rxd_7[0]~q ;
wire \rxd_7[0]~_wirecell_combout ;
wire \rxd_0[4]~q ;
wire \rxd_1[4]~q ;
wire \rxd_0[7]~q ;
wire \rxd_1[7]~q ;
wire \rxd_0[6]~q ;
wire \rxd_1[6]~q ;
wire \rxd_0[5]~q ;
wire \rxd_1[5]~q ;
wire \rxd_0[3]~q ;
wire \rxd_1[3]~q ;
wire \rxd_0[2]~q ;
wire \rxd_1[2]~q ;
wire \rxd_0[1]~q ;
wire \rxd_1[1]~q ;
wire \always8~1_combout ;
wire \no_align_err_reg~0_combout ;
wire \no_align_err_reg~q ;
wire \always8~0_combout ;
wire \always8~2_combout ;
wire \no_align_err~q ;
wire \ok_sfd~q ;
wire \ok_sfd_p~5_combout ;
wire \ok_sfd_p[0]~q ;
wire \ok_sfd_p~4_combout ;
wire \ok_sfd_p[1]~q ;
wire \ok_sfd_p~3_combout ;
wire \ok_sfd_p[2]~q ;
wire \ok_sfd_p~2_combout ;
wire \ok_sfd_p[3]~q ;
wire \ok_sfd_p~1_combout ;
wire \ok_sfd_p[4]~q ;
wire \ok_sfd_p~0_combout ;
wire \ok_sfd_p[5]~q ;
wire \ok_sfd_p[6]~q ;
wire \rxd_2[3]~q ;
wire \rxd_3[3]~q ;
wire \rxd_4[3]~q ;
wire \rxd_5[3]~q ;
wire \rxd_6[3]~q ;
wire \rxd_7[3]~q ;
wire \rxd_8[3]~q ;
wire \rxd_2[7]~q ;
wire \rxd_3[7]~q ;
wire \rxd_4[7]~q ;
wire \rxd_5[7]~q ;
wire \rxd_6[7]~q ;
wire \rxd_7[7]~q ;
wire \rxd_8[7]~q ;
wire \rxd_2[2]~q ;
wire \rxd_3[2]~q ;
wire \rxd_4[2]~q ;
wire \rxd_5[2]~q ;
wire \rxd_2[1]~q ;
wire \rxd_3[1]~q ;
wire \rxd_4[1]~q ;
wire \rxd_5[1]~q ;
wire \rxd_6[1]~q ;
wire \rxd_6[2]~q ;
wire \always10~2_combout ;
wire \rxd_2[4]~q ;
wire \rxd_3[4]~q ;
wire \rxd_4[4]~q ;
wire \rxd_5[4]~q ;
wire \rxd_2[5]~q ;
wire \rxd_3[5]~q ;
wire \rxd_4[5]~q ;
wire \rxd_5[5]~q ;
wire \rxd_2[6]~q ;
wire \rxd_3[6]~q ;
wire \rxd_4[6]~q ;
wire \rxd_5[6]~q ;
wire \always10~3_combout ;
wire \rxd_6[4]~q ;
wire \rxd_6[5]~q ;
wire \rxd_6[6]~q ;
wire \always10~4_combout ;
wire \always10~6_combout ;
wire \rxd_7[1]~q ;
wire \rxd_8[0]~q ;
wire \rxd_8[1]~q ;
wire \rxd_7[2]~q ;
wire \rxd_7[4]~q ;
wire \rxd_7[5]~q ;
wire \rxd_7[6]~q ;
wire \always10~0_combout ;
wire \rxd_8[2]~q ;
wire \rxd_8[4]~q ;
wire \rxd_8[5]~q ;
wire \rxd_8[6]~q ;
wire \always10~1_combout ;
wire \always10~7_combout ;
wire \always10~8_combout ;
wire \always10~9_combout ;
wire \always10~10_combout ;
wire \always10~11_combout ;
wire \always10~12_combout ;
wire \unicast_mac~q ;
wire \always10~5_combout ;
wire \unicast_add~q ;
wire \WideAnd0~0_combout ;
wire \WideAnd0~combout ;
wire \broad_sub[0]~q ;
wire \broad_sub[1]~q ;
wire \broad_sub[2]~q ;
wire \broad_sub[3]~q ;
wire \broad_sub[4]~q ;
wire \broad_sub[5]~q ;
wire \always9~0_combout ;
wire \always9~1_combout ;
wire \broad_add~q ;
wire \ok_sfd_p[7]~q ;
wire \always10~14_combout ;
wire \multicast_en[0]~q ;
wire \multicast_en[1]~q ;
wire \always10~13_combout ;
wire \dest_add_ok[0]~q ;
wire \dest_add_ok[1]~q ;
wire \dest_add_ok[2]~q ;
wire \dest_add_ok[3]~q ;
wire \dest_add_ok[4]~q ;
wire \dest_add_ok[5]~q ;
wire \dest_add_ok[6]~q ;
wire \dest_add_ok[7]~q ;
wire \dest_add_ok[8]~q ;
wire \dest_add_ok[9]~q ;
wire \user_length[0]~0_combout ;
wire \user_length[0]~q ;
wire \rxd_8[2]~_wirecell_combout ;
wire \user_length[10]~q ;
wire \rxd_7[1]~_wirecell_combout ;
wire \user_length[1]~q ;
wire \rxd_7[2]~_wirecell_combout ;
wire \user_length[2]~q ;
wire \rxd_7[3]~_wirecell_combout ;
wire \user_length[3]~q ;
wire \rxd_7[4]~_wirecell_combout ;
wire \user_length[4]~q ;
wire \rxd_7[5]~_wirecell_combout ;
wire \user_length[5]~q ;
wire \always15~1_combout ;
wire \rxd_7[6]~_wirecell_combout ;
wire \user_length[6]~q ;
wire \rxd_7[7]~_wirecell_combout ;
wire \user_length[7]~q ;
wire \rxd_8[0]~_wirecell_combout ;
wire \user_length[8]~q ;
wire \rxd_8[1]~_wirecell_combout ;
wire \user_length[9]~q ;
wire \user_p_lgth_inf_46_reg~1_combout ;
wire \rxd_8[3]~_wirecell_combout ;
wire \user_length[11]~q ;
wire \rxd_8[4]~_wirecell_combout ;
wire \user_length[12]~q ;
wire \rxd_8[5]~_wirecell_combout ;
wire \user_length[13]~q ;
wire \rxd_8[6]~_wirecell_combout ;
wire \user_length[14]~q ;
wire \rxd_8[7]~_wirecell_combout ;
wire \user_length[15]~q ;
wire \user_p_lgth_inf_46_reg~0_combout ;
wire \user_length_invalid~0_combout ;
wire \user_length_invalid~q ;
wire \user_p_lgth_inf_46_reg~3_combout ;
wire \user_p_lgth_inf_46_reg[0]~q ;
wire \Add0~1_sumout ;
wire \cnt_end[0]~q ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \cnt_end[1]~q ;
wire \Equal7~0_combout ;
wire \Add0~6 ;
wire \Add0~13_sumout ;
wire \cnt_end[2]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \cnt_end[3]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \cnt_end[4]~q ;
wire \Add0~22 ;
wire \Add0~9_sumout ;
wire \cnt_end[5]~q ;
wire \Equal7~1_combout ;
wire \always13~0_combout ;
wire \always13~1_combout ;
wire \cnt_end_64_user_reg[0]~q ;
wire \cnt_end_64_user_reg[1]~q ;
wire \cnt_end_64_user_reg[2]~q ;
wire \cnt_end_64_user_reg[3]~q ;
wire \cnt_end_64_user_reg[4]~q ;
wire \cnt_end_64_user_reg[5]~q ;
wire \cnt_end_64_user_reg[6]~q ;
wire \cnt_end_64_user_reg[7]~q ;
wire \cnt_end_64_user_reg[8]~q ;
wire \cnt_end_64_user_reg[9]~q ;
wire \cnt_end_64_user_reg[10]~q ;
wire \cnt_end_64_user_reg[11]~q ;
wire \cnt_end_64_user_reg[12]~q ;
wire \cnt_end_64_user_reg[13]~q ;
wire \cnt_end_64_user_reg[14]~q ;
wire \rx_en_s[25]~q ;
wire \dest_add_ok[10]~q ;
wire \dest_add_ok[11]~q ;
wire \dest_add_ok[12]~q ;
wire \dest_pause_add_ok~0_combout ;
wire \dest_pause_add_ok~q ;
wire \always14~3_combout ;
wire \always14~4_combout ;
wire \pause_type~q ;
wire \always14~5_combout ;
wire \pause_opcode~q ;
wire \always14~1_combout ;
wire \cmd_frm[0]~q ;
wire \user_frm~0_combout ;
wire \user_frm~q ;
wire \cmd_frm[1]~q ;
wire \always14~2_combout ;
wire \frm_type_ok_s[0]~q ;
wire \always15~7_combout ;
wire \cnt_wait~q ;
wire \always15~5_combout ;
wire \cnt_res~q ;
wire \always15~6_combout ;
wire \cnt_inc~q ;
wire \Add2~45_sumout ;
wire \crc_vld[1]~q ;
wire \crc_vld[2]~q ;
wire \crc_vld[3]~q ;
wire \crc_vld[4]~q ;
wire \crc_vld[5]~q ;
wire \always15~3_combout ;
wire \adder[0]~q ;
wire \Add2~46 ;
wire \Add2~49_sumout ;
wire \adder[1]~q ;
wire \Add2~50 ;
wire \Add2~53_sumout ;
wire \adder[2]~q ;
wire \Add2~54 ;
wire \Add2~57_sumout ;
wire \adder[3]~q ;
wire \Add2~58 ;
wire \Add2~61_sumout ;
wire \adder[4]~q ;
wire \Add2~62 ;
wire \Add2~41_sumout ;
wire \adder[5]~q ;
wire \Add2~42 ;
wire \Add2~37_sumout ;
wire \adder[6]~q ;
wire \Add2~38 ;
wire \Add2~33_sumout ;
wire \adder[7]~q ;
wire \Add2~34 ;
wire \Add2~29_sumout ;
wire \adder[8]~q ;
wire \Add2~30 ;
wire \Add2~1_sumout ;
wire \adder[9]~q ;
wire \Add2~2 ;
wire \Add2~25_sumout ;
wire \adder[10]~q ;
wire \Add2~26 ;
wire \Add2~5_sumout ;
wire \adder[11]~q ;
wire \Add2~6 ;
wire \Add2~17_sumout ;
wire \adder[12]~q ;
wire \Add2~18 ;
wire \Add2~21_sumout ;
wire \adder[13]~q ;
wire \Add2~22 ;
wire \Add2~13_sumout ;
wire \adder[14]~q ;
wire \Add2~14 ;
wire \Add2~9_sumout ;
wire \adder[15]~q ;
wire \always15~0_combout ;
wire \LessThan3~0_combout ;
wire \LessThan3~1_combout ;
wire \inf_64~q ;
wire \always15~4_combout ;
wire \frm_max_eq[3]~q ;
wire \Equal14~0_combout ;
wire \frm_max_eq[2]~q ;
wire \Equal13~0_combout ;
wire \frm_max_eq[1]~q ;
wire \Equal12~0_combout ;
wire \frm_max_eq[0]~q ;
wire \Equal16~0_combout ;
wire \sup_frm_maxv~q ;
wire \always15~2_combout ;
wire \frm_lgth_err_reg[0]~q ;
wire \frm_lgth_err_reg[1]~q ;
wire \end_wr_fifo~0_combout ;
wire \end_wr_fifo~1_combout ;
wire \end_wr_fifo~q ;
wire \ok_sfd_discard~0_combout ;
wire \ok_sfd_discard~q ;
wire \ok_sfd_discard_p[0]~q ;
wire \ok_sfd_discard_p[1]~q ;
wire \ok_sfd_discard_p[2]~q ;
wire \ok_sfd_discard_p[3]~q ;
wire \ok_sfd_discard_p[4]~q ;
wire \ok_sfd_discard_p[5]~q ;
wire \ok_sfd_discard_p[6]~q ;
wire \ok_sfd_discard_p[7]~q ;
wire \ok_sfd_discard_p[8]~q ;
wire \ok_sfd_discard_p[9]~q ;
wire \ok_sfd_discard_p[10]~q ;
wire \ok_sfd_discard_p[11]~q ;
wire \ok_sfd_discard_p[12]~q ;
wire \ok_sfd_discard_p[13]~q ;
wire \ok_sfd_discard_p[14]~q ;
wire \ok_sfd_discard_p[15]~q ;
wire \ok_sfd_discard_p[16]~q ;
wire \ok_sfd_discard_p[17]~q ;
wire \ok_sfd_discard_p[18]~q ;
wire \ok_sfd_discard_p[19]~q ;
wire \ok_sfd_discard_p[20]~q ;
wire \ok_sfd_discard_p[21]~q ;
wire \always14~0_combout ;
wire \frm_to_write~q ;
wire \always20~3_combout ;
wire \start_wr_fifo~q ;
wire \always20~4_combout ;
wire \fifo_wr_wait~q ;
wire \always20~5_combout ;
wire \fifo_wr~q ;
wire \user_p_lgth_inf_46_reg~2_combout ;
wire \user_p_lgth_inf_46_reg[1]~q ;
wire \always20~8_combout ;
wire \stat_wr~q ;
wire \always20~7_combout ;
wire \stat_wr_wait~q ;
wire \rx_stat_wren_s~0_combout ;
wire \rx_stat_wren_s[0]~q ;
wire \rx_stat_wren_s[1]~q ;
wire \rx_stat_wren_s[2]~q ;
wire \rx_stat_wren_s[3]~q ;
wire \rx_stat_wren_s[4]~q ;
wire \rx_stat_wren_s[5]~q ;
wire \rx_stat_wren_s[6]~q ;
wire \rx_stat_wren_s[7]~q ;
wire \rx_stat_wren_s[8]~q ;
wire \rx_stat_wren_s[9]~q ;
wire \rx_stat_wren_s[10]~q ;
wire \rx_stat_wren_s[11]~q ;
wire \current_frame~0_combout ;
wire \current_frame~q ;
wire \sleep_mode_ena~0_combout ;
wire \sleep_mode_ena~q ;
wire \rx_stat_wren~0_combout ;
wire \payload_length[0]~1_combout ;
wire \payload_length[0]~0_combout ;
wire \payload_length[1]~2_combout ;
wire \payload_length[2]~3_combout ;
wire \payload_length[3]~4_combout ;
wire \payload_length[4]~5_combout ;
wire \payload_length[5]~6_combout ;
wire \payload_length[6]~7_combout ;
wire \payload_length[7]~8_combout ;
wire \payload_length[8]~9_combout ;
wire \payload_length[9]~10_combout ;
wire \payload_length[10]~11_combout ;
wire \payload_length[11]~12_combout ;
wire \payload_length[12]~13_combout ;
wire \payload_length[13]~14_combout ;
wire \payload_length[14]~15_combout ;
wire \payload_length[15]~16_combout ;
wire \always20~0_combout ;
wire \always20~1_combout ;
wire \gm_rx_col_reg[0]~q ;
wire \gm_rx_col_reg[1]~q ;
wire \gm_rx_col_reg[2]~q ;
wire \gm_rx_col_reg[3]~q ;
wire \col_int~0_combout ;
wire \col_int~q ;
wire \col_reg[0]~q ;
wire \col_reg[1]~q ;
wire \col_reg[2]~q ;
wire \col_reg[3]~q ;
wire \col_reg[4]~q ;
wire \col_reg[5]~q ;
wire \col_reg[6]~q ;
wire \col_reg[7]~q ;
wire \col_reg[8]~q ;
wire \col_reg[9]~q ;
wire \col_reg[10]~q ;
wire \col_reg[11]~q ;
wire \col_reg[12]~q ;
wire \col_reg[13]~q ;
wire \col_reg[14]~q ;
wire \col_reg[15]~q ;
wire \col_reg[16]~q ;
wire \col_reg[17]~q ;
wire \col_reg[18]~q ;
wire \col_reg[19]~q ;
wire \col_reg[20]~q ;
wire \col_reg[21]~q ;
wire \col_reg[22]~q ;
wire \col_reg[23]~q ;
wire \col_reg[24]~q ;
wire \col_reg[25]~q ;
wire \col_reg[26]~q ;
wire \col_reg[27]~q ;
wire \col_reg[28]~q ;
wire \col_reg[29]~q ;
wire \col_reg[30]~q ;
wire \rx_stat_data_s~0_combout ;
wire \Equal17~0_combout ;
wire \Equal17~1_combout ;
wire \Equal17~2_combout ;
wire \Equal17~3_combout ;
wire \Equal17~4_combout ;
wire \frm_length_error~0_combout ;
wire \frm_length_error~1_combout ;
wire \frm_length_error~2_combout ;
wire \frm_length_error~q ;
wire \frm_lgth_err_s_reg~0_combout ;
wire \frm_lgth_err_s_reg~q ;
wire \rx_stat_data_s~1_combout ;
wire \crc_ok[1]~q ;
wire \crc_ok[2]~q ;
wire \crc_ok[3]~q ;
wire \crc_ok[4]~q ;
wire \rx_stat_data_s~2_combout ;
wire \rx_a_full_s~0_combout ;
wire \rx_a_full_s~q ;
wire \rx_stat_data_s~3_combout ;
wire \rx_err_s~0_combout ;
wire \rx_err_s[0]~q ;
wire \rx_err_s[1]~q ;
wire \rx_err_s[2]~q ;
wire \rx_err_s[3]~q ;
wire \rx_err_s[4]~q ;
wire \rx_err_s[5]~q ;
wire \rx_err_s[6]~q ;
wire \rx_err_s[7]~q ;
wire \rx_err_s[8]~q ;
wire \rx_err_s[9]~q ;
wire \rx_err_s[10]~q ;
wire \rx_err_s[11]~q ;
wire \rx_err_s[12]~q ;
wire \rx_err_s[13]~q ;
wire \rx_err_s[14]~q ;
wire \rx_err_s[15]~q ;
wire \rx_err_s[16]~q ;
wire \rx_err_s[17]~q ;
wire \rx_err_s[18]~q ;
wire \rx_err_s[19]~q ;
wire \rx_err_s[20]~q ;
wire \rx_err_s[21]~q ;
wire \rx_err_s[22]~q ;
wire \rx_err_s[23]~q ;
wire \rx_err_latched_temp~0_combout ;
wire \rx_err_latched_temp~q ;
wire \frm_type_ok_s[1]~q ;
wire \frm_ok~0_combout ;
wire \frm_ok~q ;
wire \rx_err_latched~0_combout ;
wire \rx_err_latched~q ;
wire \rx_stat_data_s~4_combout ;
wire \always20~2_combout ;
wire \always10~15_combout ;
wire \unicast_add_reg[0]~q ;
wire \unicast_add_reg[1]~q ;
wire \unicast_add_reg[2]~q ;
wire \unicast_add_reg[3]~q ;
wire \unicast_add_reg[4]~q ;
wire \unicast_add_reg[5]~q ;
wire \unicast_add_reg[6]~q ;
wire \unicast_add_reg[7]~q ;
wire \unicast_add_reg[8]~q ;
wire \unicast_add_reg[9]~q ;
wire \unicast_add_reg[10]~q ;
wire \unicast_add_reg[11]~q ;
wire \unicast_add_reg[12]~q ;
wire \unicast_add_reg[13]~q ;
wire \unicast_add_reg[14]~q ;
wire \unicast_add_reg[15]~q ;
wire \unicast_add_reg[16]~q ;
wire \broad_add_reg~0_combout ;
wire \broad_add_reg~q ;
wire \multicast_add_reg[0]~q ;
wire \multicast_add_reg[1]~q ;
wire \multicast_add_reg[2]~q ;
wire \multicast_add_reg[3]~q ;
wire \multicast_add_reg[4]~q ;
wire \multicast_add_reg[5]~q ;
wire \multicast_add_reg[6]~q ;
wire \multicast_add_reg[7]~q ;
wire \multicast_add_reg[8]~q ;
wire \multicast_add_reg[9]~q ;
wire \multicast_add_reg[10]~q ;
wire \multicast_add_reg[11]~q ;
wire \multicast_add_reg[12]~q ;
wire \multicast_add_reg[13]~q ;
wire \multicast_add_reg[14]~q ;
wire \rx_mcast~0_combout ;
wire \rx_mcast~1_combout ;
wire \always20~6_combout ;
wire \cmd_rcv~0_combout ;
wire \always25~0_combout ;
wire \always25~1_combout ;
wire \always25~2_combout ;
wire \always25~3_combout ;
wire \always25~4_combout ;
wire \always25~5_combout ;
wire \always25~6_combout ;
wire \always25~7_combout ;
wire \rxd_25[3]~q ;
wire \rxd_25[2]~q ;
wire \rxd_25[1]~q ;
wire \rxd_25[0]~q ;
wire \rxd_25[7]~q ;
wire \rxd_25[6]~q ;
wire \rxd_25[5]~q ;
wire \rxd_25[4]~q ;


IoTOctopus_QSYS_altera_tse_crc328checker U_CRC(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.rxclk_ena(rxclk_ena),
	.eof_dly_2(\U_CRC|eof_dly[2]~q ),
	.frm_type_ok_s_0(\frm_type_ok_s[0]~q ),
	.crc_ok1(\U_CRC|crc_ok~q ),
	.rxd_25_3(\rxd_25[3]~q ),
	.rxd_25_2(\rxd_25[2]~q ),
	.rxd_25_1(\rxd_25[1]~q ),
	.rxd_25_0(\rxd_25[0]~q ),
	.rxd_25_7(\rxd_25[7]~q ),
	.rxd_25_6(\rxd_25[6]~q ),
	.rxd_25_5(\rxd_25[5]~q ),
	.rxd_25_4(\rxd_25[4]~q ),
	.eof(\eof_crc~0_combout ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_127 U_SYNC_PAD_ENA(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_PAD_ENA|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_118 U_SYNC_13(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.dreg_11(\U_SYNC_13|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_116 U_SYNC_11(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_11|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_altshifttaps U_SHIFTTAPS(
	.ram_block5a4(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout ),
	.ram_block5a5(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ),
	.ram_block5a6(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6~portbdataout ),
	.ram_block5a7(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7~portbdataout ),
	.ram_block5a0(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ),
	.ram_block5a1(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ),
	.ram_block5a2(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout ),
	.ram_block5a3(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ),
	.rxclk_ena(rxclk_ena),
	.rxd_8_0(\rxd_8[0]~q ),
	.rxd_8_1(\rxd_8[1]~q ),
	.rxd_8_2(\rxd_8[2]~q ),
	.rxd_8_3(\rxd_8[3]~q ),
	.rxd_8_4(\rxd_8[4]~q ),
	.rxd_8_5(\rxd_8[5]~q ),
	.rxd_8_6(\rxd_8[6]~q ),
	.rxd_8_7(\rxd_8[7]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_115 U_SYNC_10(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.ethernet_mode(ethernet_mode),
	.dreg_1(\U_SYNC_10|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_126 U_SYNC_9(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_9|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_124 U_SYNC_7(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_7|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_123 U_SYNC_6(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_121 U_SYNC_4(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_120 U_SYNC_3(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_3|std_sync_no_cut|dreg[1]~q ),
	.sleep_ena(sleep_ena),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_119 U_SYNC_2(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_114 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.mac_rx_clock_connection_clk(mac_rx_clock_connection_clk));

cyclonev_lcell_comb \eof_crc~0 (
	.dataa(!\rx_en_s[24]~q ),
	.datab(!\rx_en_s[23]~q ),
	.datac(!\frm_ok~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eof_crc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eof_crc~0 .extended_lut = "off";
defparam \eof_crc~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \eof_crc~0 .shared_arith = "off";

dffeas rx_stat_wren(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_stat_wren1),
	.prn(vcc));
defparam rx_stat_wren.is_wysiwyg = "true";
defparam rx_stat_wren.power_up = "low";

dffeas \payload_length[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_0),
	.prn(vcc));
defparam \payload_length[0] .is_wysiwyg = "true";
defparam \payload_length[0] .power_up = "low";

dffeas \payload_length[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_1),
	.prn(vcc));
defparam \payload_length[1] .is_wysiwyg = "true";
defparam \payload_length[1] .power_up = "low";

dffeas \payload_length[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_2),
	.prn(vcc));
defparam \payload_length[2] .is_wysiwyg = "true";
defparam \payload_length[2] .power_up = "low";

dffeas \payload_length[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_3),
	.prn(vcc));
defparam \payload_length[3] .is_wysiwyg = "true";
defparam \payload_length[3] .power_up = "low";

dffeas \payload_length[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[4]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_4),
	.prn(vcc));
defparam \payload_length[4] .is_wysiwyg = "true";
defparam \payload_length[4] .power_up = "low";

dffeas \payload_length[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[5]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_5),
	.prn(vcc));
defparam \payload_length[5] .is_wysiwyg = "true";
defparam \payload_length[5] .power_up = "low";

dffeas \payload_length[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[6]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_6),
	.prn(vcc));
defparam \payload_length[6] .is_wysiwyg = "true";
defparam \payload_length[6] .power_up = "low";

dffeas \payload_length[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[7]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_7),
	.prn(vcc));
defparam \payload_length[7] .is_wysiwyg = "true";
defparam \payload_length[7] .power_up = "low";

dffeas \payload_length[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[8]~9_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_8),
	.prn(vcc));
defparam \payload_length[8] .is_wysiwyg = "true";
defparam \payload_length[8] .power_up = "low";

dffeas \payload_length[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[9]~10_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_9),
	.prn(vcc));
defparam \payload_length[9] .is_wysiwyg = "true";
defparam \payload_length[9] .power_up = "low";

dffeas \payload_length[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[10]~11_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_10),
	.prn(vcc));
defparam \payload_length[10] .is_wysiwyg = "true";
defparam \payload_length[10] .power_up = "low";

dffeas \payload_length[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[11]~12_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_11),
	.prn(vcc));
defparam \payload_length[11] .is_wysiwyg = "true";
defparam \payload_length[11] .power_up = "low";

dffeas \payload_length[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[12]~13_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_12),
	.prn(vcc));
defparam \payload_length[12] .is_wysiwyg = "true";
defparam \payload_length[12] .power_up = "low";

dffeas \payload_length[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[13]~14_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_13),
	.prn(vcc));
defparam \payload_length[13] .is_wysiwyg = "true";
defparam \payload_length[13] .power_up = "low";

dffeas \payload_length[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[14]~15_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_14),
	.prn(vcc));
defparam \payload_length[14] .is_wysiwyg = "true";
defparam \payload_length[14] .power_up = "low";

dffeas \payload_length[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\payload_length[15]~16_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\payload_length[0]~0_combout ),
	.q(payload_length_15),
	.prn(vcc));
defparam \payload_length[15] .is_wysiwyg = "true";
defparam \payload_length[15] .power_up = "low";

dffeas rx_wren_int(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_wren_int1),
	.prn(vcc));
defparam rx_wren_int.is_wysiwyg = "true";
defparam rx_wren_int.power_up = "low";

dffeas rx_eop_int(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_eop_int1),
	.prn(vcc));
defparam rx_eop_int.is_wysiwyg = "true";
defparam rx_eop_int.power_up = "low";

dffeas \rx_stat_data_s[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_data_s~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_stat_data_s_5),
	.prn(vcc));
defparam \rx_stat_data_s[5] .is_wysiwyg = "true";
defparam \rx_stat_data_s[5] .power_up = "low";

dffeas \rx_stat_data_s[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_data_s~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_stat_data_s_0),
	.prn(vcc));
defparam \rx_stat_data_s[0] .is_wysiwyg = "true";
defparam \rx_stat_data_s[0] .power_up = "low";

dffeas \rx_stat_data_s[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_data_s~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_stat_data_s_1),
	.prn(vcc));
defparam \rx_stat_data_s[1] .is_wysiwyg = "true";
defparam \rx_stat_data_s[1] .power_up = "low";

dffeas \rx_stat_data_s[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_data_s~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_stat_data_s_2),
	.prn(vcc));
defparam \rx_stat_data_s[2] .is_wysiwyg = "true";
defparam \rx_stat_data_s[2] .power_up = "low";

dffeas \rx_stat_data_s[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_data_s~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_stat_data_s_3),
	.prn(vcc));
defparam \rx_stat_data_s[3] .is_wysiwyg = "true";
defparam \rx_stat_data_s[3] .power_up = "low";

dffeas rx_sop_int(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_sop_int1),
	.prn(vcc));
defparam rx_sop_int.is_wysiwyg = "true";
defparam rx_sop_int.power_up = "low";

dffeas rx_ucast(
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[16]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_ucast1),
	.prn(vcc));
defparam rx_ucast.is_wysiwyg = "true";
defparam rx_ucast.power_up = "low";

dffeas rx_mcast(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_mcast~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_mcast1),
	.prn(vcc));
defparam rx_mcast.is_wysiwyg = "true";
defparam rx_mcast.power_up = "low";

dffeas rx_bcast(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_mcast~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_bcast1),
	.prn(vcc));
defparam rx_bcast.is_wysiwyg = "true";
defparam rx_bcast.power_up = "low";

dffeas rx_data_val(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_val1),
	.prn(vcc));
defparam rx_data_val.is_wysiwyg = "true";
defparam rx_data_val.power_up = "low";

dffeas magic_pkt_ena(
	.clk(mac_rx_clock_connection_clk),
	.d(\cmd_rcv~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(magic_pkt_ena1),
	.prn(vcc));
defparam magic_pkt_ena.is_wysiwyg = "true";
defparam magic_pkt_ena.power_up = "low";

dffeas rx_done_reg(
	.clk(mac_rx_clock_connection_clk),
	.d(\always25~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rx_done_reg1),
	.prn(vcc));
defparam rx_done_reg.is_wysiwyg = "true";
defparam rx_done_reg.power_up = "low";

dffeas \rx_data_int[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_3),
	.prn(vcc));
defparam \rx_data_int[3] .is_wysiwyg = "true";
defparam \rx_data_int[3] .power_up = "low";

dffeas \rx_data_int[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_2),
	.prn(vcc));
defparam \rx_data_int[2] .is_wysiwyg = "true";
defparam \rx_data_int[2] .power_up = "low";

dffeas \rx_data_int[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_1),
	.prn(vcc));
defparam \rx_data_int[1] .is_wysiwyg = "true";
defparam \rx_data_int[1] .power_up = "low";

dffeas \rx_data_int[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_0),
	.prn(vcc));
defparam \rx_data_int[0] .is_wysiwyg = "true";
defparam \rx_data_int[0] .power_up = "low";

dffeas \rx_data_int[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_7),
	.prn(vcc));
defparam \rx_data_int[7] .is_wysiwyg = "true";
defparam \rx_data_int[7] .power_up = "low";

dffeas \rx_data_int[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_6),
	.prn(vcc));
defparam \rx_data_int[6] .is_wysiwyg = "true";
defparam \rx_data_int[6] .power_up = "low";

dffeas \rx_data_int[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_5),
	.prn(vcc));
defparam \rx_data_int[5] .is_wysiwyg = "true";
defparam \rx_data_int[5] .power_up = "low";

dffeas \rx_data_int[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_25[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(rx_data_int_4),
	.prn(vcc));
defparam \rx_data_int[4] .is_wysiwyg = "true";
defparam \rx_data_int[4] .power_up = "low";

cyclonev_lcell_comb \enable_rx_reg3~0 (
	.dataa(!\enable_rx_reg3~q ),
	.datab(!en),
	.datac(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\enable_rx_reg3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \enable_rx_reg3~0 .extended_lut = "off";
defparam \enable_rx_reg3~0 .lut_mask = 64'h4747474747474747;
defparam \enable_rx_reg3~0 .shared_arith = "off";

dffeas enable_rx_reg3(
	.clk(mac_rx_clock_connection_clk),
	.d(\enable_rx_reg3~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\enable_rx_reg3~q ),
	.prn(vcc));
defparam enable_rx_reg3.is_wysiwyg = "true";
defparam enable_rx_reg3.power_up = "low";

cyclonev_lcell_comb \rx_en_s~0 (
	.dataa(!\enable_rx_reg3~q ),
	.datab(!en),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_en_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_en_s~0 .extended_lut = "off";
defparam \rx_en_s~0 .lut_mask = 64'h7777777777777777;
defparam \rx_en_s~0 .shared_arith = "off";

dffeas \rx_en_s[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[0]~q ),
	.prn(vcc));
defparam \rx_en_s[0] .is_wysiwyg = "true";
defparam \rx_en_s[0] .power_up = "low";

dffeas \rx_en_s[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[1]~q ),
	.prn(vcc));
defparam \rx_en_s[1] .is_wysiwyg = "true";
defparam \rx_en_s[1] .power_up = "low";

dffeas \rx_en_s[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[2]~q ),
	.prn(vcc));
defparam \rx_en_s[2] .is_wysiwyg = "true";
defparam \rx_en_s[2] .power_up = "low";

dffeas \rx_en_s[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[3]~q ),
	.prn(vcc));
defparam \rx_en_s[3] .is_wysiwyg = "true";
defparam \rx_en_s[3] .power_up = "low";

dffeas \rx_en_s[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[4]~q ),
	.prn(vcc));
defparam \rx_en_s[4] .is_wysiwyg = "true";
defparam \rx_en_s[4] .power_up = "low";

dffeas \rx_en_s[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[5]~q ),
	.prn(vcc));
defparam \rx_en_s[5] .is_wysiwyg = "true";
defparam \rx_en_s[5] .power_up = "low";

dffeas \rx_en_s[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[6]~q ),
	.prn(vcc));
defparam \rx_en_s[6] .is_wysiwyg = "true";
defparam \rx_en_s[6] .power_up = "low";

dffeas \rx_en_s[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[7]~q ),
	.prn(vcc));
defparam \rx_en_s[7] .is_wysiwyg = "true";
defparam \rx_en_s[7] .power_up = "low";

dffeas \rx_en_s[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[8]~q ),
	.prn(vcc));
defparam \rx_en_s[8] .is_wysiwyg = "true";
defparam \rx_en_s[8] .power_up = "low";

dffeas \rx_en_s[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[9]~q ),
	.prn(vcc));
defparam \rx_en_s[9] .is_wysiwyg = "true";
defparam \rx_en_s[9] .power_up = "low";

dffeas \rx_en_s[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[10]~q ),
	.prn(vcc));
defparam \rx_en_s[10] .is_wysiwyg = "true";
defparam \rx_en_s[10] .power_up = "low";

dffeas \rx_en_s[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[11]~q ),
	.prn(vcc));
defparam \rx_en_s[11] .is_wysiwyg = "true";
defparam \rx_en_s[11] .power_up = "low";

dffeas \rx_en_s[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[12]~q ),
	.prn(vcc));
defparam \rx_en_s[12] .is_wysiwyg = "true";
defparam \rx_en_s[12] .power_up = "low";

dffeas \rx_en_s[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[13]~q ),
	.prn(vcc));
defparam \rx_en_s[13] .is_wysiwyg = "true";
defparam \rx_en_s[13] .power_up = "low";

dffeas \rx_en_s[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[14]~q ),
	.prn(vcc));
defparam \rx_en_s[14] .is_wysiwyg = "true";
defparam \rx_en_s[14] .power_up = "low";

dffeas \rx_en_s[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[14]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[15]~q ),
	.prn(vcc));
defparam \rx_en_s[15] .is_wysiwyg = "true";
defparam \rx_en_s[15] .power_up = "low";

dffeas \rx_en_s[16] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[15]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[16]~q ),
	.prn(vcc));
defparam \rx_en_s[16] .is_wysiwyg = "true";
defparam \rx_en_s[16] .power_up = "low";

dffeas \rx_en_s[17] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[16]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[17]~q ),
	.prn(vcc));
defparam \rx_en_s[17] .is_wysiwyg = "true";
defparam \rx_en_s[17] .power_up = "low";

dffeas \rx_en_s[18] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[17]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[18]~q ),
	.prn(vcc));
defparam \rx_en_s[18] .is_wysiwyg = "true";
defparam \rx_en_s[18] .power_up = "low";

dffeas \rx_en_s[19] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[18]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[19]~q ),
	.prn(vcc));
defparam \rx_en_s[19] .is_wysiwyg = "true";
defparam \rx_en_s[19] .power_up = "low";

dffeas \rx_en_s[20] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[19]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[20]~q ),
	.prn(vcc));
defparam \rx_en_s[20] .is_wysiwyg = "true";
defparam \rx_en_s[20] .power_up = "low";

dffeas \rx_en_s[21] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[20]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[21]~q ),
	.prn(vcc));
defparam \rx_en_s[21] .is_wysiwyg = "true";
defparam \rx_en_s[21] .power_up = "low";

dffeas \rx_en_s[22] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[21]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[22]~q ),
	.prn(vcc));
defparam \rx_en_s[22] .is_wysiwyg = "true";
defparam \rx_en_s[22] .power_up = "low";

dffeas \rx_en_s[23] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[22]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[23]~q ),
	.prn(vcc));
defparam \rx_en_s[23] .is_wysiwyg = "true";
defparam \rx_en_s[23] .power_up = "low";

dffeas \rx_en_s[24] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[23]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[24]~q ),
	.prn(vcc));
defparam \rx_en_s[24] .is_wysiwyg = "true";
defparam \rx_en_s[24] .power_up = "low";

dffeas \rxd_0[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[0]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[0]~q ),
	.prn(vcc));
defparam \rxd_0[0] .is_wysiwyg = "true";
defparam \rxd_0[0] .power_up = "low";

dffeas \rxd_1[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[0]~q ),
	.prn(vcc));
defparam \rxd_1[0] .is_wysiwyg = "true";
defparam \rxd_1[0] .power_up = "low";

dffeas \rxd_2[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[0]~q ),
	.prn(vcc));
defparam \rxd_2[0] .is_wysiwyg = "true";
defparam \rxd_2[0] .power_up = "low";

dffeas \rxd_3[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[0]~q ),
	.prn(vcc));
defparam \rxd_3[0] .is_wysiwyg = "true";
defparam \rxd_3[0] .power_up = "low";

dffeas \rxd_4[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[0]~q ),
	.prn(vcc));
defparam \rxd_4[0] .is_wysiwyg = "true";
defparam \rxd_4[0] .power_up = "low";

dffeas \rxd_5[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[0]~q ),
	.prn(vcc));
defparam \rxd_5[0] .is_wysiwyg = "true";
defparam \rxd_5[0] .power_up = "low";

dffeas \rxd_6[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[0]~q ),
	.prn(vcc));
defparam \rxd_6[0] .is_wysiwyg = "true";
defparam \rxd_6[0] .power_up = "low";

dffeas \rxd_7[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[0]~q ),
	.prn(vcc));
defparam \rxd_7[0] .is_wysiwyg = "true";
defparam \rxd_7[0] .power_up = "low";

cyclonev_lcell_comb \rxd_7[0]~_wirecell (
	.dataa(!\rxd_7[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[0]~_wirecell .extended_lut = "off";
defparam \rxd_7[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[0]~_wirecell .shared_arith = "off";

dffeas \rxd_0[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[4]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[4]~q ),
	.prn(vcc));
defparam \rxd_0[4] .is_wysiwyg = "true";
defparam \rxd_0[4] .power_up = "low";

dffeas \rxd_1[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[4]~q ),
	.prn(vcc));
defparam \rxd_1[4] .is_wysiwyg = "true";
defparam \rxd_1[4] .power_up = "low";

dffeas \rxd_0[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[7]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[7]~q ),
	.prn(vcc));
defparam \rxd_0[7] .is_wysiwyg = "true";
defparam \rxd_0[7] .power_up = "low";

dffeas \rxd_1[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[7]~q ),
	.prn(vcc));
defparam \rxd_1[7] .is_wysiwyg = "true";
defparam \rxd_1[7] .power_up = "low";

dffeas \rxd_0[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[6]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[6]~q ),
	.prn(vcc));
defparam \rxd_0[6] .is_wysiwyg = "true";
defparam \rxd_0[6] .power_up = "low";

dffeas \rxd_1[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[6]~q ),
	.prn(vcc));
defparam \rxd_1[6] .is_wysiwyg = "true";
defparam \rxd_1[6] .power_up = "low";

dffeas \rxd_0[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[5]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[5]~q ),
	.prn(vcc));
defparam \rxd_0[5] .is_wysiwyg = "true";
defparam \rxd_0[5] .power_up = "low";

dffeas \rxd_1[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[5]~q ),
	.prn(vcc));
defparam \rxd_1[5] .is_wysiwyg = "true";
defparam \rxd_1[5] .power_up = "low";

dffeas \rxd_0[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[3]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[3]~q ),
	.prn(vcc));
defparam \rxd_0[3] .is_wysiwyg = "true";
defparam \rxd_0[3] .power_up = "low";

dffeas \rxd_1[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[3]~q ),
	.prn(vcc));
defparam \rxd_1[3] .is_wysiwyg = "true";
defparam \rxd_1[3] .power_up = "low";

dffeas \rxd_0[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[2]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[2]~q ),
	.prn(vcc));
defparam \rxd_0[2] .is_wysiwyg = "true";
defparam \rxd_0[2] .power_up = "low";

dffeas \rxd_1[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[2]~q ),
	.prn(vcc));
defparam \rxd_1[2] .is_wysiwyg = "true";
defparam \rxd_1[2] .power_up = "low";

dffeas \rxd_0[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(rx_d[1]),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_0[1]~q ),
	.prn(vcc));
defparam \rxd_0[1] .is_wysiwyg = "true";
defparam \rxd_0[1] .power_up = "low";

dffeas \rxd_1[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_0[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\enable_rx_reg3~q ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_1[1]~q ),
	.prn(vcc));
defparam \rxd_1[1] .is_wysiwyg = "true";
defparam \rxd_1[1] .power_up = "low";

cyclonev_lcell_comb \always8~1 (
	.dataa(!\rxd_1[3]~q ),
	.datab(!\rxd_1[2]~q ),
	.datac(!\rxd_1[1]~q ),
	.datad(!\rxd_1[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always8~1 .extended_lut = "off";
defparam \always8~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \always8~1 .shared_arith = "off";

cyclonev_lcell_comb \no_align_err_reg~0 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rxd_1[4]~q ),
	.datac(!\no_align_err_reg~q ),
	.datad(!\always8~0_combout ),
	.datae(!\always8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\no_align_err_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \no_align_err_reg~0 .extended_lut = "off";
defparam \no_align_err_reg~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \no_align_err_reg~0 .shared_arith = "off";

dffeas no_align_err_reg(
	.clk(mac_rx_clock_connection_clk),
	.d(\no_align_err_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\no_align_err_reg~q ),
	.prn(vcc));
defparam no_align_err_reg.is_wysiwyg = "true";
defparam no_align_err_reg.power_up = "low";

cyclonev_lcell_comb \always8~0 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rxd_1[7]~q ),
	.datac(!\rxd_1[6]~q ),
	.datad(!\rxd_1[5]~q ),
	.datae(!\no_align_err_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always8~0 .extended_lut = "off";
defparam \always8~0 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \always8~0 .shared_arith = "off";

cyclonev_lcell_comb \always8~2 (
	.dataa(!\rxd_1[4]~q ),
	.datab(!\always8~0_combout ),
	.datac(!\always8~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always8~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always8~2 .extended_lut = "off";
defparam \always8~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always8~2 .shared_arith = "off";

dffeas no_align_err(
	.clk(mac_rx_clock_connection_clk),
	.d(\always8~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\no_align_err~q ),
	.prn(vcc));
defparam no_align_err.is_wysiwyg = "true";
defparam no_align_err.power_up = "low";

dffeas ok_sfd(
	.clk(mac_rx_clock_connection_clk),
	.d(\no_align_err~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd~q ),
	.prn(vcc));
defparam ok_sfd.is_wysiwyg = "true";
defparam ok_sfd.power_up = "low";

cyclonev_lcell_comb \ok_sfd_p~5 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rx_en_s[0]~q ),
	.datac(!\ok_sfd~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_p~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_p~5 .extended_lut = "off";
defparam \ok_sfd_p~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ok_sfd_p~5 .shared_arith = "off";

dffeas \ok_sfd_p[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[0]~q ),
	.prn(vcc));
defparam \ok_sfd_p[0] .is_wysiwyg = "true";
defparam \ok_sfd_p[0] .power_up = "low";

cyclonev_lcell_comb \ok_sfd_p~4 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rx_en_s[0]~q ),
	.datac(!\ok_sfd_p[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_p~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_p~4 .extended_lut = "off";
defparam \ok_sfd_p~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ok_sfd_p~4 .shared_arith = "off";

dffeas \ok_sfd_p[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[1]~q ),
	.prn(vcc));
defparam \ok_sfd_p[1] .is_wysiwyg = "true";
defparam \ok_sfd_p[1] .power_up = "low";

cyclonev_lcell_comb \ok_sfd_p~3 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rx_en_s[0]~q ),
	.datac(!\ok_sfd_p[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_p~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_p~3 .extended_lut = "off";
defparam \ok_sfd_p~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ok_sfd_p~3 .shared_arith = "off";

dffeas \ok_sfd_p[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[2]~q ),
	.prn(vcc));
defparam \ok_sfd_p[2] .is_wysiwyg = "true";
defparam \ok_sfd_p[2] .power_up = "low";

cyclonev_lcell_comb \ok_sfd_p~2 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rx_en_s[0]~q ),
	.datac(!\ok_sfd_p[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_p~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_p~2 .extended_lut = "off";
defparam \ok_sfd_p~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ok_sfd_p~2 .shared_arith = "off";

dffeas \ok_sfd_p[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[3]~q ),
	.prn(vcc));
defparam \ok_sfd_p[3] .is_wysiwyg = "true";
defparam \ok_sfd_p[3] .power_up = "low";

cyclonev_lcell_comb \ok_sfd_p~1 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rx_en_s[0]~q ),
	.datac(!\ok_sfd_p[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_p~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_p~1 .extended_lut = "off";
defparam \ok_sfd_p~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ok_sfd_p~1 .shared_arith = "off";

dffeas \ok_sfd_p[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[4]~q ),
	.prn(vcc));
defparam \ok_sfd_p[4] .is_wysiwyg = "true";
defparam \ok_sfd_p[4] .power_up = "low";

cyclonev_lcell_comb \ok_sfd_p~0 (
	.dataa(!\rx_en_s[1]~q ),
	.datab(!\rx_en_s[0]~q ),
	.datac(!\ok_sfd_p[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_p~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_p~0 .extended_lut = "off";
defparam \ok_sfd_p~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ok_sfd_p~0 .shared_arith = "off";

dffeas \ok_sfd_p[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[5]~q ),
	.prn(vcc));
defparam \ok_sfd_p[5] .is_wysiwyg = "true";
defparam \ok_sfd_p[5] .power_up = "low";

dffeas \ok_sfd_p[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[6]~q ),
	.prn(vcc));
defparam \ok_sfd_p[6] .is_wysiwyg = "true";
defparam \ok_sfd_p[6] .power_up = "low";

dffeas \rxd_2[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[3]~q ),
	.prn(vcc));
defparam \rxd_2[3] .is_wysiwyg = "true";
defparam \rxd_2[3] .power_up = "low";

dffeas \rxd_3[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[3]~q ),
	.prn(vcc));
defparam \rxd_3[3] .is_wysiwyg = "true";
defparam \rxd_3[3] .power_up = "low";

dffeas \rxd_4[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[3]~q ),
	.prn(vcc));
defparam \rxd_4[3] .is_wysiwyg = "true";
defparam \rxd_4[3] .power_up = "low";

dffeas \rxd_5[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[3]~q ),
	.prn(vcc));
defparam \rxd_5[3] .is_wysiwyg = "true";
defparam \rxd_5[3] .power_up = "low";

dffeas \rxd_6[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[3]~q ),
	.prn(vcc));
defparam \rxd_6[3] .is_wysiwyg = "true";
defparam \rxd_6[3] .power_up = "low";

dffeas \rxd_7[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[3]~q ),
	.prn(vcc));
defparam \rxd_7[3] .is_wysiwyg = "true";
defparam \rxd_7[3] .power_up = "low";

dffeas \rxd_8[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[3]~q ),
	.prn(vcc));
defparam \rxd_8[3] .is_wysiwyg = "true";
defparam \rxd_8[3] .power_up = "low";

dffeas \rxd_2[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[7]~q ),
	.prn(vcc));
defparam \rxd_2[7] .is_wysiwyg = "true";
defparam \rxd_2[7] .power_up = "low";

dffeas \rxd_3[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[7]~q ),
	.prn(vcc));
defparam \rxd_3[7] .is_wysiwyg = "true";
defparam \rxd_3[7] .power_up = "low";

dffeas \rxd_4[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[7]~q ),
	.prn(vcc));
defparam \rxd_4[7] .is_wysiwyg = "true";
defparam \rxd_4[7] .power_up = "low";

dffeas \rxd_5[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[7]~q ),
	.prn(vcc));
defparam \rxd_5[7] .is_wysiwyg = "true";
defparam \rxd_5[7] .power_up = "low";

dffeas \rxd_6[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[7]~q ),
	.prn(vcc));
defparam \rxd_6[7] .is_wysiwyg = "true";
defparam \rxd_6[7] .power_up = "low";

dffeas \rxd_7[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[7]~q ),
	.prn(vcc));
defparam \rxd_7[7] .is_wysiwyg = "true";
defparam \rxd_7[7] .power_up = "low";

dffeas \rxd_8[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[7]~q ),
	.prn(vcc));
defparam \rxd_8[7] .is_wysiwyg = "true";
defparam \rxd_8[7] .power_up = "low";

dffeas \rxd_2[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[2]~q ),
	.prn(vcc));
defparam \rxd_2[2] .is_wysiwyg = "true";
defparam \rxd_2[2] .power_up = "low";

dffeas \rxd_3[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[2]~q ),
	.prn(vcc));
defparam \rxd_3[2] .is_wysiwyg = "true";
defparam \rxd_3[2] .power_up = "low";

dffeas \rxd_4[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[2]~q ),
	.prn(vcc));
defparam \rxd_4[2] .is_wysiwyg = "true";
defparam \rxd_4[2] .power_up = "low";

dffeas \rxd_5[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[2]~q ),
	.prn(vcc));
defparam \rxd_5[2] .is_wysiwyg = "true";
defparam \rxd_5[2] .power_up = "low";

dffeas \rxd_2[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[1]~q ),
	.prn(vcc));
defparam \rxd_2[1] .is_wysiwyg = "true";
defparam \rxd_2[1] .power_up = "low";

dffeas \rxd_3[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[1]~q ),
	.prn(vcc));
defparam \rxd_3[1] .is_wysiwyg = "true";
defparam \rxd_3[1] .power_up = "low";

dffeas \rxd_4[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[1]~q ),
	.prn(vcc));
defparam \rxd_4[1] .is_wysiwyg = "true";
defparam \rxd_4[1] .power_up = "low";

dffeas \rxd_5[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[1]~q ),
	.prn(vcc));
defparam \rxd_5[1] .is_wysiwyg = "true";
defparam \rxd_5[1] .power_up = "low";

dffeas \rxd_6[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[1]~q ),
	.prn(vcc));
defparam \rxd_6[1] .is_wysiwyg = "true";
defparam \rxd_6[1] .power_up = "low";

dffeas \rxd_6[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[2]~q ),
	.prn(vcc));
defparam \rxd_6[2] .is_wysiwyg = "true";
defparam \rxd_6[2] .power_up = "low";

cyclonev_lcell_comb \always10~2 (
	.dataa(!\rxd_6[0]~q ),
	.datab(!\rxd_6[1]~q ),
	.datac(!\rxd_6[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~2 .extended_lut = "off";
defparam \always10~2 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \always10~2 .shared_arith = "off";

dffeas \rxd_2[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[4]~q ),
	.prn(vcc));
defparam \rxd_2[4] .is_wysiwyg = "true";
defparam \rxd_2[4] .power_up = "low";

dffeas \rxd_3[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[4]~q ),
	.prn(vcc));
defparam \rxd_3[4] .is_wysiwyg = "true";
defparam \rxd_3[4] .power_up = "low";

dffeas \rxd_4[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[4]~q ),
	.prn(vcc));
defparam \rxd_4[4] .is_wysiwyg = "true";
defparam \rxd_4[4] .power_up = "low";

dffeas \rxd_5[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[4]~q ),
	.prn(vcc));
defparam \rxd_5[4] .is_wysiwyg = "true";
defparam \rxd_5[4] .power_up = "low";

dffeas \rxd_2[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[5]~q ),
	.prn(vcc));
defparam \rxd_2[5] .is_wysiwyg = "true";
defparam \rxd_2[5] .power_up = "low";

dffeas \rxd_3[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[5]~q ),
	.prn(vcc));
defparam \rxd_3[5] .is_wysiwyg = "true";
defparam \rxd_3[5] .power_up = "low";

dffeas \rxd_4[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[5]~q ),
	.prn(vcc));
defparam \rxd_4[5] .is_wysiwyg = "true";
defparam \rxd_4[5] .power_up = "low";

dffeas \rxd_5[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[5]~q ),
	.prn(vcc));
defparam \rxd_5[5] .is_wysiwyg = "true";
defparam \rxd_5[5] .power_up = "low";

dffeas \rxd_2[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_1[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_2[6]~q ),
	.prn(vcc));
defparam \rxd_2[6] .is_wysiwyg = "true";
defparam \rxd_2[6] .power_up = "low";

dffeas \rxd_3[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_2[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_3[6]~q ),
	.prn(vcc));
defparam \rxd_3[6] .is_wysiwyg = "true";
defparam \rxd_3[6] .power_up = "low";

dffeas \rxd_4[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_3[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_4[6]~q ),
	.prn(vcc));
defparam \rxd_4[6] .is_wysiwyg = "true";
defparam \rxd_4[6] .power_up = "low";

dffeas \rxd_5[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_4[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_5[6]~q ),
	.prn(vcc));
defparam \rxd_5[6] .is_wysiwyg = "true";
defparam \rxd_5[6] .power_up = "low";

cyclonev_lcell_comb \always10~3 (
	.dataa(!\rxd_5[3]~q ),
	.datab(!\rxd_5[4]~q ),
	.datac(!\rxd_5[5]~q ),
	.datad(!\rxd_5[6]~q ),
	.datae(!\rxd_5[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~3 .extended_lut = "off";
defparam \always10~3 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~3 .shared_arith = "off";

dffeas \rxd_6[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[4]~q ),
	.prn(vcc));
defparam \rxd_6[4] .is_wysiwyg = "true";
defparam \rxd_6[4] .power_up = "low";

dffeas \rxd_6[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[5]~q ),
	.prn(vcc));
defparam \rxd_6[5] .is_wysiwyg = "true";
defparam \rxd_6[5] .power_up = "low";

dffeas \rxd_6[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_5[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_6[6]~q ),
	.prn(vcc));
defparam \rxd_6[6] .is_wysiwyg = "true";
defparam \rxd_6[6] .power_up = "low";

cyclonev_lcell_comb \always10~4 (
	.dataa(!\rxd_6[4]~q ),
	.datab(!\rxd_6[5]~q ),
	.datac(!\rxd_6[6]~q ),
	.datad(!\rxd_6[7]~q ),
	.datae(!\rxd_5[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~4 .extended_lut = "off";
defparam \always10~4 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~4 .shared_arith = "off";

cyclonev_lcell_comb \always10~6 (
	.dataa(!\rxd_6[3]~q ),
	.datab(!\rxd_5[2]~q ),
	.datac(!\always10~2_combout ),
	.datad(!\always10~3_combout ),
	.datae(!\always10~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~6 .extended_lut = "off";
defparam \always10~6 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \always10~6 .shared_arith = "off";

dffeas \rxd_7[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[1]~q ),
	.prn(vcc));
defparam \rxd_7[1] .is_wysiwyg = "true";
defparam \rxd_7[1] .power_up = "low";

dffeas \rxd_8[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[0]~q ),
	.prn(vcc));
defparam \rxd_8[0] .is_wysiwyg = "true";
defparam \rxd_8[0] .power_up = "low";

dffeas \rxd_8[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[1]~q ),
	.prn(vcc));
defparam \rxd_8[1] .is_wysiwyg = "true";
defparam \rxd_8[1] .power_up = "low";

dffeas \rxd_7[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[2]~q ),
	.prn(vcc));
defparam \rxd_7[2] .is_wysiwyg = "true";
defparam \rxd_7[2] .power_up = "low";

dffeas \rxd_7[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[4]~q ),
	.prn(vcc));
defparam \rxd_7[4] .is_wysiwyg = "true";
defparam \rxd_7[4] .power_up = "low";

dffeas \rxd_7[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[5]~q ),
	.prn(vcc));
defparam \rxd_7[5] .is_wysiwyg = "true";
defparam \rxd_7[5] .power_up = "low";

dffeas \rxd_7[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_6[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_7[6]~q ),
	.prn(vcc));
defparam \rxd_7[6] .is_wysiwyg = "true";
defparam \rxd_7[6] .power_up = "low";

cyclonev_lcell_comb \always10~0 (
	.dataa(!\rxd_7[2]~q ),
	.datab(!\rxd_7[4]~q ),
	.datac(!\rxd_7[5]~q ),
	.datad(!\rxd_7[6]~q ),
	.datae(!\rxd_7[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~0 .shared_arith = "off";

dffeas \rxd_8[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[2]~q ),
	.prn(vcc));
defparam \rxd_8[2] .is_wysiwyg = "true";
defparam \rxd_8[2] .power_up = "low";

dffeas \rxd_8[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[4]~q ),
	.prn(vcc));
defparam \rxd_8[4] .is_wysiwyg = "true";
defparam \rxd_8[4] .power_up = "low";

dffeas \rxd_8[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[5]~q ),
	.prn(vcc));
defparam \rxd_8[5] .is_wysiwyg = "true";
defparam \rxd_8[5] .power_up = "low";

dffeas \rxd_8[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rxd_7[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_8[6]~q ),
	.prn(vcc));
defparam \rxd_8[6] .is_wysiwyg = "true";
defparam \rxd_8[6] .power_up = "low";

cyclonev_lcell_comb \always10~1 (
	.dataa(!\rxd_7[0]~q ),
	.datab(!\rxd_8[2]~q ),
	.datac(!\rxd_8[4]~q ),
	.datad(!\rxd_8[5]~q ),
	.datae(!\rxd_8[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "off";
defparam \always10~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \always10~7 (
	.dataa(!\rxd_7[1]~q ),
	.datab(!\rxd_8[0]~q ),
	.datac(!\rxd_8[1]~q ),
	.datad(!\always10~0_combout ),
	.datae(!\always10~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~7 .extended_lut = "off";
defparam \always10~7 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \always10~7 .shared_arith = "off";

cyclonev_lcell_comb \always10~8 (
	.dataa(!\rxd_3[7]~q ),
	.datab(!\rxd_3[6]~q ),
	.datac(!\rxd_3[5]~q ),
	.datad(!\rxd_3[4]~q ),
	.datae(!\rxd_3[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~8 .extended_lut = "off";
defparam \always10~8 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~8 .shared_arith = "off";

cyclonev_lcell_comb \always10~9 (
	.dataa(!\rxd_3[1]~q ),
	.datab(!\rxd_3[0]~q ),
	.datac(!\rxd_4[5]~q ),
	.datad(!\rxd_4[6]~q ),
	.datae(!\rxd_4[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~9 .extended_lut = "off";
defparam \always10~9 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~9 .shared_arith = "off";

cyclonev_lcell_comb \always10~10 (
	.dataa(!\rxd_5[0]~q ),
	.datab(!\rxd_4[0]~q ),
	.datac(!\rxd_4[1]~q ),
	.datad(!\rxd_4[2]~q ),
	.datae(!\rxd_4[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~10 .extended_lut = "off";
defparam \always10~10 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always10~10 .shared_arith = "off";

cyclonev_lcell_comb \always10~11 (
	.dataa(!\rxd_7[3]~q ),
	.datab(!\rxd_3[2]~q ),
	.datac(!\rxd_4[4]~q ),
	.datad(!\always10~8_combout ),
	.datae(!\always10~9_combout ),
	.dataf(!\always10~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~11 .extended_lut = "off";
defparam \always10~11 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \always10~11 .shared_arith = "off";

cyclonev_lcell_comb \always10~12 (
	.dataa(!\rxd_8[3]~q ),
	.datab(!\rxd_8[7]~q ),
	.datac(!\always10~6_combout ),
	.datad(!\always10~7_combout ),
	.datae(!\always10~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~12 .extended_lut = "off";
defparam \always10~12 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \always10~12 .shared_arith = "off";

dffeas unicast_mac(
	.clk(mac_rx_clock_connection_clk),
	.d(\always10~12_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_mac~q ),
	.prn(vcc));
defparam unicast_mac.is_wysiwyg = "true";
defparam unicast_mac.power_up = "low";

cyclonev_lcell_comb \always10~5 (
	.dataa(!\ok_sfd_p[6]~q ),
	.datab(!\unicast_mac~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~5 .extended_lut = "off";
defparam \always10~5 .lut_mask = 64'h7777777777777777;
defparam \always10~5 .shared_arith = "off";

dffeas unicast_add(
	.clk(mac_rx_clock_connection_clk),
	.d(\always10~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add~q ),
	.prn(vcc));
defparam unicast_add.is_wysiwyg = "true";
defparam unicast_add.power_up = "low";

cyclonev_lcell_comb \WideAnd0~0 (
	.dataa(!\rxd_3[7]~q ),
	.datab(!\rxd_3[6]~q ),
	.datac(!\rxd_3[5]~q ),
	.datad(!\rxd_3[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideAnd0~0 .extended_lut = "off";
defparam \WideAnd0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \WideAnd0~0 .shared_arith = "off";

cyclonev_lcell_comb WideAnd0(
	.dataa(!\rxd_3[3]~q ),
	.datab(!\rxd_3[2]~q ),
	.datac(!\rxd_3[1]~q ),
	.datad(!\rxd_3[0]~q ),
	.datae(!\WideAnd0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideAnd0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam WideAnd0.extended_lut = "off";
defparam WideAnd0.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam WideAnd0.shared_arith = "off";

dffeas \broad_sub[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\WideAnd0~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_sub[0]~q ),
	.prn(vcc));
defparam \broad_sub[0] .is_wysiwyg = "true";
defparam \broad_sub[0] .power_up = "low";

dffeas \broad_sub[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\broad_sub[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_sub[1]~q ),
	.prn(vcc));
defparam \broad_sub[1] .is_wysiwyg = "true";
defparam \broad_sub[1] .power_up = "low";

dffeas \broad_sub[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\broad_sub[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_sub[2]~q ),
	.prn(vcc));
defparam \broad_sub[2] .is_wysiwyg = "true";
defparam \broad_sub[2] .power_up = "low";

dffeas \broad_sub[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\broad_sub[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_sub[3]~q ),
	.prn(vcc));
defparam \broad_sub[3] .is_wysiwyg = "true";
defparam \broad_sub[3] .power_up = "low";

dffeas \broad_sub[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\broad_sub[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_sub[4]~q ),
	.prn(vcc));
defparam \broad_sub[4] .is_wysiwyg = "true";
defparam \broad_sub[4] .power_up = "low";

dffeas \broad_sub[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\broad_sub[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_sub[5]~q ),
	.prn(vcc));
defparam \broad_sub[5] .is_wysiwyg = "true";
defparam \broad_sub[5] .power_up = "low";

cyclonev_lcell_comb \always9~0 (
	.dataa(!\broad_sub[5]~q ),
	.datab(!\broad_sub[4]~q ),
	.datac(!\broad_sub[3]~q ),
	.datad(!\broad_sub[2]~q ),
	.datae(!\broad_sub[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \always9~0 .shared_arith = "off";

cyclonev_lcell_comb \always9~1 (
	.dataa(!\broad_sub[0]~q ),
	.datab(!\ok_sfd_p[6]~q ),
	.datac(!\always9~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~1 .extended_lut = "off";
defparam \always9~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always9~1 .shared_arith = "off";

dffeas broad_add(
	.clk(mac_rx_clock_connection_clk),
	.d(\always9~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_add~q ),
	.prn(vcc));
defparam broad_add.is_wysiwyg = "true";
defparam broad_add.power_up = "low";

dffeas \ok_sfd_p[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_p[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_p[7]~q ),
	.prn(vcc));
defparam \ok_sfd_p[7] .is_wysiwyg = "true";
defparam \ok_sfd_p[7] .power_up = "low";

cyclonev_lcell_comb \always10~14 (
	.dataa(!\rxd_8[0]~q ),
	.datab(!\ok_sfd_p[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~14 .extended_lut = "off";
defparam \always10~14 .lut_mask = 64'h7777777777777777;
defparam \always10~14 .shared_arith = "off";

dffeas \multicast_en[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always10~14_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_en[0]~q ),
	.prn(vcc));
defparam \multicast_en[0] .is_wysiwyg = "true";
defparam \multicast_en[0] .power_up = "low";

dffeas \multicast_en[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_en[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_en[1]~q ),
	.prn(vcc));
defparam \multicast_en[1] .is_wysiwyg = "true";
defparam \multicast_en[1] .power_up = "low";

cyclonev_lcell_comb \always10~13 (
	.dataa(!\unicast_add~q ),
	.datab(!\broad_add~q ),
	.datac(!\ok_sfd_p[7]~q ),
	.datad(!\U_SYNC_9|std_sync_no_cut|dreg[1]~q ),
	.datae(!\multicast_en[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~13 .extended_lut = "off";
defparam \always10~13 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \always10~13 .shared_arith = "off";

dffeas \dest_add_ok[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always10~13_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[0]~q ),
	.prn(vcc));
defparam \dest_add_ok[0] .is_wysiwyg = "true";
defparam \dest_add_ok[0] .power_up = "low";

dffeas \dest_add_ok[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[1]~q ),
	.prn(vcc));
defparam \dest_add_ok[1] .is_wysiwyg = "true";
defparam \dest_add_ok[1] .power_up = "low";

dffeas \dest_add_ok[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[2]~q ),
	.prn(vcc));
defparam \dest_add_ok[2] .is_wysiwyg = "true";
defparam \dest_add_ok[2] .power_up = "low";

dffeas \dest_add_ok[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[3]~q ),
	.prn(vcc));
defparam \dest_add_ok[3] .is_wysiwyg = "true";
defparam \dest_add_ok[3] .power_up = "low";

dffeas \dest_add_ok[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[4]~q ),
	.prn(vcc));
defparam \dest_add_ok[4] .is_wysiwyg = "true";
defparam \dest_add_ok[4] .power_up = "low";

dffeas \dest_add_ok[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[5]~q ),
	.prn(vcc));
defparam \dest_add_ok[5] .is_wysiwyg = "true";
defparam \dest_add_ok[5] .power_up = "low";

dffeas \dest_add_ok[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[6]~q ),
	.prn(vcc));
defparam \dest_add_ok[6] .is_wysiwyg = "true";
defparam \dest_add_ok[6] .power_up = "low";

dffeas \dest_add_ok[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[7]~q ),
	.prn(vcc));
defparam \dest_add_ok[7] .is_wysiwyg = "true";
defparam \dest_add_ok[7] .power_up = "low";

dffeas \dest_add_ok[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[8]~q ),
	.prn(vcc));
defparam \dest_add_ok[8] .is_wysiwyg = "true";
defparam \dest_add_ok[8] .power_up = "low";

dffeas \dest_add_ok[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[9]~q ),
	.prn(vcc));
defparam \dest_add_ok[9] .is_wysiwyg = "true";
defparam \dest_add_ok[9] .power_up = "low";

cyclonev_lcell_comb \user_length[0]~0 (
	.dataa(!rxclk_ena),
	.datab(!\dest_add_ok[9]~q ),
	.datac(!\rx_en_s[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_length[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_length[0]~0 .extended_lut = "off";
defparam \user_length[0]~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \user_length[0]~0 .shared_arith = "off";

dffeas \user_length[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[0]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[0]~q ),
	.prn(vcc));
defparam \user_length[0] .is_wysiwyg = "true";
defparam \user_length[0] .power_up = "low";

cyclonev_lcell_comb \rxd_8[2]~_wirecell (
	.dataa(!\rxd_8[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[2]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[2]~_wirecell .extended_lut = "off";
defparam \rxd_8[2]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[2]~_wirecell .shared_arith = "off";

dffeas \user_length[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[2]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[10]~q ),
	.prn(vcc));
defparam \user_length[10] .is_wysiwyg = "true";
defparam \user_length[10] .power_up = "low";

cyclonev_lcell_comb \rxd_7[1]~_wirecell (
	.dataa(!\rxd_7[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[1]~_wirecell .extended_lut = "off";
defparam \rxd_7[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[1]~_wirecell .shared_arith = "off";

dffeas \user_length[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[1]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[1]~q ),
	.prn(vcc));
defparam \user_length[1] .is_wysiwyg = "true";
defparam \user_length[1] .power_up = "low";

cyclonev_lcell_comb \rxd_7[2]~_wirecell (
	.dataa(!\rxd_7[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[2]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[2]~_wirecell .extended_lut = "off";
defparam \rxd_7[2]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[2]~_wirecell .shared_arith = "off";

dffeas \user_length[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[2]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[2]~q ),
	.prn(vcc));
defparam \user_length[2] .is_wysiwyg = "true";
defparam \user_length[2] .power_up = "low";

cyclonev_lcell_comb \rxd_7[3]~_wirecell (
	.dataa(!\rxd_7[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[3]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[3]~_wirecell .extended_lut = "off";
defparam \rxd_7[3]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[3]~_wirecell .shared_arith = "off";

dffeas \user_length[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[3]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[3]~q ),
	.prn(vcc));
defparam \user_length[3] .is_wysiwyg = "true";
defparam \user_length[3] .power_up = "low";

cyclonev_lcell_comb \rxd_7[4]~_wirecell (
	.dataa(!\rxd_7[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[4]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[4]~_wirecell .extended_lut = "off";
defparam \rxd_7[4]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[4]~_wirecell .shared_arith = "off";

dffeas \user_length[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[4]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[4]~q ),
	.prn(vcc));
defparam \user_length[4] .is_wysiwyg = "true";
defparam \user_length[4] .power_up = "low";

cyclonev_lcell_comb \rxd_7[5]~_wirecell (
	.dataa(!\rxd_7[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[5]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[5]~_wirecell .extended_lut = "off";
defparam \rxd_7[5]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[5]~_wirecell .shared_arith = "off";

dffeas \user_length[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[5]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[5]~q ),
	.prn(vcc));
defparam \user_length[5] .is_wysiwyg = "true";
defparam \user_length[5] .power_up = "low";

cyclonev_lcell_comb \always15~1 (
	.dataa(!\user_length[1]~q ),
	.datab(!\user_length[2]~q ),
	.datac(!\user_length[3]~q ),
	.datad(!\user_length[4]~q ),
	.datae(!\user_length[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~1 .extended_lut = "off";
defparam \always15~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always15~1 .shared_arith = "off";

cyclonev_lcell_comb \rxd_7[6]~_wirecell (
	.dataa(!\rxd_7[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[6]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[6]~_wirecell .extended_lut = "off";
defparam \rxd_7[6]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[6]~_wirecell .shared_arith = "off";

dffeas \user_length[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[6]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[6]~q ),
	.prn(vcc));
defparam \user_length[6] .is_wysiwyg = "true";
defparam \user_length[6] .power_up = "low";

cyclonev_lcell_comb \rxd_7[7]~_wirecell (
	.dataa(!\rxd_7[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_7[7]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_7[7]~_wirecell .extended_lut = "off";
defparam \rxd_7[7]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_7[7]~_wirecell .shared_arith = "off";

dffeas \user_length[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_7[7]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[7]~q ),
	.prn(vcc));
defparam \user_length[7] .is_wysiwyg = "true";
defparam \user_length[7] .power_up = "low";

cyclonev_lcell_comb \rxd_8[0]~_wirecell (
	.dataa(!\rxd_8[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[0]~_wirecell .extended_lut = "off";
defparam \rxd_8[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[0]~_wirecell .shared_arith = "off";

dffeas \user_length[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[0]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[8]~q ),
	.prn(vcc));
defparam \user_length[8] .is_wysiwyg = "true";
defparam \user_length[8] .power_up = "low";

cyclonev_lcell_comb \rxd_8[1]~_wirecell (
	.dataa(!\rxd_8[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[1]~_wirecell .extended_lut = "off";
defparam \rxd_8[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[1]~_wirecell .shared_arith = "off";

dffeas \user_length[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[1]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[9]~q ),
	.prn(vcc));
defparam \user_length[9] .is_wysiwyg = "true";
defparam \user_length[9] .power_up = "low";

cyclonev_lcell_comb \user_p_lgth_inf_46_reg~1 (
	.dataa(!\user_length[6]~q ),
	.datab(!\user_length[7]~q ),
	.datac(!\user_length[8]~q ),
	.datad(!\user_length[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_p_lgth_inf_46_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_p_lgth_inf_46_reg~1 .extended_lut = "off";
defparam \user_p_lgth_inf_46_reg~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \user_p_lgth_inf_46_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \rxd_8[3]~_wirecell (
	.dataa(!\rxd_8[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[3]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[3]~_wirecell .extended_lut = "off";
defparam \rxd_8[3]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[3]~_wirecell .shared_arith = "off";

dffeas \user_length[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[3]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[11]~q ),
	.prn(vcc));
defparam \user_length[11] .is_wysiwyg = "true";
defparam \user_length[11] .power_up = "low";

cyclonev_lcell_comb \rxd_8[4]~_wirecell (
	.dataa(!\rxd_8[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[4]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[4]~_wirecell .extended_lut = "off";
defparam \rxd_8[4]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[4]~_wirecell .shared_arith = "off";

dffeas \user_length[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[4]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[12]~q ),
	.prn(vcc));
defparam \user_length[12] .is_wysiwyg = "true";
defparam \user_length[12] .power_up = "low";

cyclonev_lcell_comb \rxd_8[5]~_wirecell (
	.dataa(!\rxd_8[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[5]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[5]~_wirecell .extended_lut = "off";
defparam \rxd_8[5]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[5]~_wirecell .shared_arith = "off";

dffeas \user_length[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[5]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[13]~q ),
	.prn(vcc));
defparam \user_length[13] .is_wysiwyg = "true";
defparam \user_length[13] .power_up = "low";

cyclonev_lcell_comb \rxd_8[6]~_wirecell (
	.dataa(!\rxd_8[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[6]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[6]~_wirecell .extended_lut = "off";
defparam \rxd_8[6]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[6]~_wirecell .shared_arith = "off";

dffeas \user_length[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[6]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[14]~q ),
	.prn(vcc));
defparam \user_length[14] .is_wysiwyg = "true";
defparam \user_length[14] .power_up = "low";

cyclonev_lcell_comb \rxd_8[7]~_wirecell (
	.dataa(!\rxd_8[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rxd_8[7]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rxd_8[7]~_wirecell .extended_lut = "off";
defparam \rxd_8[7]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \rxd_8[7]~_wirecell .shared_arith = "off";

dffeas \user_length[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rxd_8[7]~_wirecell_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(\user_length[0]~0_combout ),
	.q(\user_length[15]~q ),
	.prn(vcc));
defparam \user_length[15] .is_wysiwyg = "true";
defparam \user_length[15] .power_up = "low";

cyclonev_lcell_comb \user_p_lgth_inf_46_reg~0 (
	.dataa(!\user_length[11]~q ),
	.datab(!\user_length[12]~q ),
	.datac(!\user_length[13]~q ),
	.datad(!\user_length[14]~q ),
	.datae(!\user_length[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_p_lgth_inf_46_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_p_lgth_inf_46_reg~0 .extended_lut = "off";
defparam \user_p_lgth_inf_46_reg~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \user_p_lgth_inf_46_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \user_length_invalid~0 (
	.dataa(!\dest_add_ok[9]~q ),
	.datab(!\rx_en_s[14]~q ),
	.datac(!\rx_en_s[7]~q ),
	.datad(!\user_length_invalid~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_length_invalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_length_invalid~0 .extended_lut = "off";
defparam \user_length_invalid~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \user_length_invalid~0 .shared_arith = "off";

dffeas user_length_invalid(
	.clk(mac_rx_clock_connection_clk),
	.d(\user_length_invalid~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\user_length_invalid~q ),
	.prn(vcc));
defparam user_length_invalid.is_wysiwyg = "true";
defparam user_length_invalid.power_up = "low";

cyclonev_lcell_comb \user_p_lgth_inf_46_reg~3 (
	.dataa(!\user_length[10]~q ),
	.datab(!\always15~1_combout ),
	.datac(!\user_p_lgth_inf_46_reg~1_combout ),
	.datad(!\user_p_lgth_inf_46_reg~0_combout ),
	.datae(!\user_length_invalid~q ),
	.dataf(!\U_SYNC_PAD_ENA|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_p_lgth_inf_46_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_p_lgth_inf_46_reg~3 .extended_lut = "off";
defparam \user_p_lgth_inf_46_reg~3 .lut_mask = 64'hFFFFDFFFFFFFFFFF;
defparam \user_p_lgth_inf_46_reg~3 .shared_arith = "off";

dffeas \user_p_lgth_inf_46_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\user_p_lgth_inf_46_reg~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\user_p_lgth_inf_46_reg[0]~q ),
	.prn(vcc));
defparam \user_p_lgth_inf_46_reg[0] .is_wysiwyg = "true";
defparam \user_p_lgth_inf_46_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt_end[0]~q ),
	.datae(gnd),
	.dataf(!\user_p_lgth_inf_46_reg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \cnt_end[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~1_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(rxclk_ena),
	.q(\cnt_end[0]~q ),
	.prn(vcc));
defparam \cnt_end[0] .is_wysiwyg = "true";
defparam \cnt_end[0] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt_end[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \cnt_end[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~5_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(rxclk_ena),
	.q(\cnt_end[1]~q ),
	.prn(vcc));
defparam \cnt_end[1] .is_wysiwyg = "true";
defparam \cnt_end[1] .power_up = "low";

cyclonev_lcell_comb \Equal7~0 (
	.dataa(!\user_length[1]~q ),
	.datab(!\cnt_end[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal7~0 .extended_lut = "off";
defparam \Equal7~0 .lut_mask = 64'h6666666666666666;
defparam \Equal7~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt_end[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \cnt_end[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~13_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(rxclk_ena),
	.q(\cnt_end[2]~q ),
	.prn(vcc));
defparam \cnt_end[2] .is_wysiwyg = "true";
defparam \cnt_end[2] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt_end[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \cnt_end[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~17_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(rxclk_ena),
	.q(\cnt_end[3]~q ),
	.prn(vcc));
defparam \cnt_end[3] .is_wysiwyg = "true";
defparam \cnt_end[3] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt_end[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \cnt_end[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~21_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(rxclk_ena),
	.q(\cnt_end[4]~q ),
	.prn(vcc));
defparam \cnt_end[4] .is_wysiwyg = "true";
defparam \cnt_end[4] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\cnt_end[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \cnt_end[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add0~9_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\dest_add_ok[9]~q ),
	.ena(rxclk_ena),
	.q(\cnt_end[5]~q ),
	.prn(vcc));
defparam \cnt_end[5] .is_wysiwyg = "true";
defparam \cnt_end[5] .power_up = "low";

cyclonev_lcell_comb \Equal7~1 (
	.dataa(!\user_length[5]~q ),
	.datab(!\cnt_end[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal7~1 .extended_lut = "off";
defparam \Equal7~1 .lut_mask = 64'h6666666666666666;
defparam \Equal7~1 .shared_arith = "off";

cyclonev_lcell_comb \always13~0 (
	.dataa(!\user_length[2]~q ),
	.datab(!\user_length[3]~q ),
	.datac(!\user_length[4]~q ),
	.datad(!\cnt_end[2]~q ),
	.datae(!\cnt_end[3]~q ),
	.dataf(!\cnt_end[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~0 .extended_lut = "off";
defparam \always13~0 .lut_mask = 64'h6996966996696996;
defparam \always13~0 .shared_arith = "off";

cyclonev_lcell_comb \always13~1 (
	.dataa(!\user_length[0]~q ),
	.datab(!\user_p_lgth_inf_46_reg[0]~q ),
	.datac(!\cnt_end[0]~q ),
	.datad(!\Equal7~0_combout ),
	.datae(!\Equal7~1_combout ),
	.dataf(!\always13~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~1 .extended_lut = "off";
defparam \always13~1 .lut_mask = 64'h7BFFFFFFFFFFFFFF;
defparam \always13~1 .shared_arith = "off";

dffeas \cnt_end_64_user_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always13~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[0]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[0] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[0] .power_up = "low";

dffeas \cnt_end_64_user_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[1]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[1] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[1] .power_up = "low";

dffeas \cnt_end_64_user_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[2]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[2] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[2] .power_up = "low";

dffeas \cnt_end_64_user_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[3]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[3] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[3] .power_up = "low";

dffeas \cnt_end_64_user_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[4]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[4] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[4] .power_up = "low";

dffeas \cnt_end_64_user_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[5]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[5] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[5] .power_up = "low";

dffeas \cnt_end_64_user_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[6]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[6] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[6] .power_up = "low";

dffeas \cnt_end_64_user_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[7]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[7] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[7] .power_up = "low";

dffeas \cnt_end_64_user_reg[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[8]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[8] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[8] .power_up = "low";

dffeas \cnt_end_64_user_reg[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[9]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[9] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[9] .power_up = "low";

dffeas \cnt_end_64_user_reg[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[10]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[10] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[10] .power_up = "low";

dffeas \cnt_end_64_user_reg[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[11]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[11] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[11] .power_up = "low";

dffeas \cnt_end_64_user_reg[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[12]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[12] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[12] .power_up = "low";

dffeas \cnt_end_64_user_reg[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[13]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[13] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[13] .power_up = "low";

dffeas \cnt_end_64_user_reg[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cnt_end_64_user_reg[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_end_64_user_reg[14]~q ),
	.prn(vcc));
defparam \cnt_end_64_user_reg[14] .is_wysiwyg = "true";
defparam \cnt_end_64_user_reg[14] .power_up = "low";

dffeas \rx_en_s[25] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_en_s[24]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_en_s[25]~q ),
	.prn(vcc));
defparam \rx_en_s[25] .is_wysiwyg = "true";
defparam \rx_en_s[25] .power_up = "low";

dffeas \dest_add_ok[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[10]~q ),
	.prn(vcc));
defparam \dest_add_ok[10] .is_wysiwyg = "true";
defparam \dest_add_ok[10] .power_up = "low";

dffeas \dest_add_ok[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[11]~q ),
	.prn(vcc));
defparam \dest_add_ok[11] .is_wysiwyg = "true";
defparam \dest_add_ok[11] .power_up = "low";

dffeas \dest_add_ok[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_add_ok[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_add_ok[12]~q ),
	.prn(vcc));
defparam \dest_add_ok[12] .is_wysiwyg = "true";
defparam \dest_add_ok[12] .power_up = "low";

cyclonev_lcell_comb \dest_pause_add_ok~0 (
	.dataa(!\dest_add_ok[11]~q ),
	.datab(!\dest_pause_add_ok~q ),
	.datac(!\unicast_add~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dest_pause_add_ok~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dest_pause_add_ok~0 .extended_lut = "off";
defparam \dest_pause_add_ok~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \dest_pause_add_ok~0 .shared_arith = "off";

dffeas dest_pause_add_ok(
	.clk(mac_rx_clock_connection_clk),
	.d(\dest_pause_add_ok~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\dest_pause_add_ok~q ),
	.prn(vcc));
defparam dest_pause_add_ok.is_wysiwyg = "true";
defparam dest_pause_add_ok.power_up = "low";

cyclonev_lcell_comb \always14~3 (
	.dataa(!\rxd_7[3]~q ),
	.datab(!\rxd_8[3]~q ),
	.datac(!\rxd_8[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~3 .extended_lut = "off";
defparam \always14~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always14~3 .shared_arith = "off";

cyclonev_lcell_comb \always14~4 (
	.dataa(!\rxd_7[1]~q ),
	.datab(!\rxd_8[0]~q ),
	.datac(!\rxd_8[1]~q ),
	.datad(!\always10~0_combout ),
	.datae(!\always10~1_combout ),
	.dataf(!\always14~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~4 .extended_lut = "off";
defparam \always14~4 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \always14~4 .shared_arith = "off";

dffeas pause_type(
	.clk(mac_rx_clock_connection_clk),
	.d(\always14~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\pause_type~q ),
	.prn(vcc));
defparam pause_type.is_wysiwyg = "true";
defparam pause_type.power_up = "low";

cyclonev_lcell_comb \always14~5 (
	.dataa(!\rxd_6[3]~q ),
	.datab(!\rxd_5[0]~q ),
	.datac(!\rxd_5[2]~q ),
	.datad(!\always10~2_combout ),
	.datae(!\always10~3_combout ),
	.dataf(!\always10~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~5 .extended_lut = "off";
defparam \always14~5 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \always14~5 .shared_arith = "off";

dffeas pause_opcode(
	.clk(mac_rx_clock_connection_clk),
	.d(\always14~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\pause_opcode~q ),
	.prn(vcc));
defparam pause_opcode.is_wysiwyg = "true";
defparam pause_opcode.power_up = "low";

cyclonev_lcell_comb \always14~1 (
	.dataa(!\dest_add_ok[10]~q ),
	.datab(!\dest_pause_add_ok~q ),
	.datac(!\pause_type~q ),
	.datad(!\pause_opcode~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~1 .extended_lut = "off";
defparam \always14~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \always14~1 .shared_arith = "off";

dffeas \cmd_frm[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always14~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cmd_frm[0]~q ),
	.prn(vcc));
defparam \cmd_frm[0] .is_wysiwyg = "true";
defparam \cmd_frm[0] .power_up = "low";

cyclonev_lcell_comb \user_frm~0 (
	.dataa(!\dest_add_ok[11]~q ),
	.datab(!\cmd_frm[0]~q ),
	.datac(!\U_SYNC_6|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_frm~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_frm~0 .extended_lut = "off";
defparam \user_frm~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \user_frm~0 .shared_arith = "off";

dffeas user_frm(
	.clk(mac_rx_clock_connection_clk),
	.d(\user_frm~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\user_frm~q ),
	.prn(vcc));
defparam user_frm.is_wysiwyg = "true";
defparam user_frm.power_up = "low";

dffeas \cmd_frm[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\cmd_frm[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cmd_frm[1]~q ),
	.prn(vcc));
defparam \cmd_frm[1] .is_wysiwyg = "true";
defparam \cmd_frm[1] .power_up = "low";

cyclonev_lcell_comb \always14~2 (
	.dataa(!\dest_add_ok[12]~q ),
	.datab(!\user_frm~q ),
	.datac(!\cmd_frm[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~2 .extended_lut = "off";
defparam \always14~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always14~2 .shared_arith = "off";

dffeas \frm_type_ok_s[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always14~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_type_ok_s[0]~q ),
	.prn(vcc));
defparam \frm_type_ok_s[0] .is_wysiwyg = "true";
defparam \frm_type_ok_s[0] .power_up = "low";

cyclonev_lcell_comb \always15~7 (
	.dataa(!\rx_en_s[24]~q ),
	.datab(!\cnt_inc~q ),
	.datac(!\frm_type_ok_s[0]~q ),
	.datad(!\cnt_wait~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~7 .extended_lut = "off";
defparam \always15~7 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \always15~7 .shared_arith = "off";

dffeas cnt_wait(
	.clk(mac_rx_clock_connection_clk),
	.d(\always15~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_wait~q ),
	.prn(vcc));
defparam cnt_wait.is_wysiwyg = "true";
defparam cnt_wait.power_up = "low";

cyclonev_lcell_comb \always15~5 (
	.dataa(!\frm_type_ok_s[0]~q ),
	.datab(!\cnt_wait~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~5 .extended_lut = "off";
defparam \always15~5 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always15~5 .shared_arith = "off";

dffeas cnt_res(
	.clk(mac_rx_clock_connection_clk),
	.d(\always15~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_res~q ),
	.prn(vcc));
defparam cnt_res.is_wysiwyg = "true";
defparam cnt_res.power_up = "low";

cyclonev_lcell_comb \always15~6 (
	.dataa(!\rx_en_s[25]~q ),
	.datab(!\cnt_inc~q ),
	.datac(!\cnt_res~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~6 .extended_lut = "off";
defparam \always15~6 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always15~6 .shared_arith = "off";

dffeas cnt_inc(
	.clk(mac_rx_clock_connection_clk),
	.d(\always15~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\cnt_inc~q ),
	.prn(vcc));
defparam cnt_inc.is_wysiwyg = "true";
defparam cnt_inc.power_up = "low";

cyclonev_lcell_comb \Add2~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[0]~q ),
	.datae(gnd),
	.dataf(!\cnt_inc~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~45_sumout ),
	.cout(\Add2~46 ),
	.shareout());
defparam \Add2~45 .extended_lut = "off";
defparam \Add2~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add2~45 .shared_arith = "off";

dffeas \crc_vld[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_CRC|eof_dly[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_vld[1]~q ),
	.prn(vcc));
defparam \crc_vld[1] .is_wysiwyg = "true";
defparam \crc_vld[1] .power_up = "low";

dffeas \crc_vld[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_vld[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_vld[2]~q ),
	.prn(vcc));
defparam \crc_vld[2] .is_wysiwyg = "true";
defparam \crc_vld[2] .power_up = "low";

dffeas \crc_vld[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_vld[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_vld[3]~q ),
	.prn(vcc));
defparam \crc_vld[3] .is_wysiwyg = "true";
defparam \crc_vld[3] .power_up = "low";

dffeas \crc_vld[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_vld[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_vld[4]~q ),
	.prn(vcc));
defparam \crc_vld[4] .is_wysiwyg = "true";
defparam \crc_vld[4] .power_up = "low";

dffeas \crc_vld[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_vld[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_vld[5]~q ),
	.prn(vcc));
defparam \crc_vld[5] .is_wysiwyg = "true";
defparam \crc_vld[5] .power_up = "low";

cyclonev_lcell_comb \always15~3 (
	.dataa(!\crc_vld[5]~q ),
	.datab(!\cnt_res~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~3 .extended_lut = "off";
defparam \always15~3 .lut_mask = 64'h7777777777777777;
defparam \always15~3 .shared_arith = "off";

dffeas \adder[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~45_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[0]~q ),
	.prn(vcc));
defparam \adder[0] .is_wysiwyg = "true";
defparam \adder[0] .power_up = "low";

cyclonev_lcell_comb \Add2~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~49_sumout ),
	.cout(\Add2~50 ),
	.shareout());
defparam \Add2~49 .extended_lut = "off";
defparam \Add2~49 .lut_mask = 64'h00000000000000FF;
defparam \Add2~49 .shared_arith = "off";

dffeas \adder[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~49_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[1]~q ),
	.prn(vcc));
defparam \adder[1] .is_wysiwyg = "true";
defparam \adder[1] .power_up = "low";

cyclonev_lcell_comb \Add2~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~53_sumout ),
	.cout(\Add2~54 ),
	.shareout());
defparam \Add2~53 .extended_lut = "off";
defparam \Add2~53 .lut_mask = 64'h00000000000000FF;
defparam \Add2~53 .shared_arith = "off";

dffeas \adder[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~53_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[2]~q ),
	.prn(vcc));
defparam \adder[2] .is_wysiwyg = "true";
defparam \adder[2] .power_up = "low";

cyclonev_lcell_comb \Add2~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~57_sumout ),
	.cout(\Add2~58 ),
	.shareout());
defparam \Add2~57 .extended_lut = "off";
defparam \Add2~57 .lut_mask = 64'h00000000000000FF;
defparam \Add2~57 .shared_arith = "off";

dffeas \adder[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~57_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[3]~q ),
	.prn(vcc));
defparam \adder[3] .is_wysiwyg = "true";
defparam \adder[3] .power_up = "low";

cyclonev_lcell_comb \Add2~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~61_sumout ),
	.cout(\Add2~62 ),
	.shareout());
defparam \Add2~61 .extended_lut = "off";
defparam \Add2~61 .lut_mask = 64'h00000000000000FF;
defparam \Add2~61 .shared_arith = "off";

dffeas \adder[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~61_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[4]~q ),
	.prn(vcc));
defparam \adder[4] .is_wysiwyg = "true";
defparam \adder[4] .power_up = "low";

cyclonev_lcell_comb \Add2~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~41_sumout ),
	.cout(\Add2~42 ),
	.shareout());
defparam \Add2~41 .extended_lut = "off";
defparam \Add2~41 .lut_mask = 64'h00000000000000FF;
defparam \Add2~41 .shared_arith = "off";

dffeas \adder[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~41_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[5]~q ),
	.prn(vcc));
defparam \adder[5] .is_wysiwyg = "true";
defparam \adder[5] .power_up = "low";

cyclonev_lcell_comb \Add2~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~37_sumout ),
	.cout(\Add2~38 ),
	.shareout());
defparam \Add2~37 .extended_lut = "off";
defparam \Add2~37 .lut_mask = 64'h00000000000000FF;
defparam \Add2~37 .shared_arith = "off";

dffeas \adder[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~37_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[6]~q ),
	.prn(vcc));
defparam \adder[6] .is_wysiwyg = "true";
defparam \adder[6] .power_up = "low";

cyclonev_lcell_comb \Add2~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~33_sumout ),
	.cout(\Add2~34 ),
	.shareout());
defparam \Add2~33 .extended_lut = "off";
defparam \Add2~33 .lut_mask = 64'h00000000000000FF;
defparam \Add2~33 .shared_arith = "off";

dffeas \adder[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~33_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[7]~q ),
	.prn(vcc));
defparam \adder[7] .is_wysiwyg = "true";
defparam \adder[7] .power_up = "low";

cyclonev_lcell_comb \Add2~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~29_sumout ),
	.cout(\Add2~30 ),
	.shareout());
defparam \Add2~29 .extended_lut = "off";
defparam \Add2~29 .lut_mask = 64'h00000000000000FF;
defparam \Add2~29 .shared_arith = "off";

dffeas \adder[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~29_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[8]~q ),
	.prn(vcc));
defparam \adder[8] .is_wysiwyg = "true";
defparam \adder[8] .power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h00000000000000FF;
defparam \Add2~1 .shared_arith = "off";

dffeas \adder[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[9]~q ),
	.prn(vcc));
defparam \adder[9] .is_wysiwyg = "true";
defparam \adder[9] .power_up = "low";

cyclonev_lcell_comb \Add2~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(\Add2~26 ),
	.shareout());
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h00000000000000FF;
defparam \Add2~25 .shared_arith = "off";

dffeas \adder[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~25_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[10]~q ),
	.prn(vcc));
defparam \adder[10] .is_wysiwyg = "true";
defparam \adder[10] .power_up = "low";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(\Add2~6 ),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h00000000000000FF;
defparam \Add2~5 .shared_arith = "off";

dffeas \adder[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[11]~q ),
	.prn(vcc));
defparam \adder[11] .is_wysiwyg = "true";
defparam \adder[11] .power_up = "low";

cyclonev_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h00000000000000FF;
defparam \Add2~17 .shared_arith = "off";

dffeas \adder[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[12]~q ),
	.prn(vcc));
defparam \adder[12] .is_wysiwyg = "true";
defparam \adder[12] .power_up = "low";

cyclonev_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h00000000000000FF;
defparam \Add2~21 .shared_arith = "off";

dffeas \adder[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~21_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[13]~q ),
	.prn(vcc));
defparam \adder[13] .is_wysiwyg = "true";
defparam \adder[13] .power_up = "low";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h00000000000000FF;
defparam \Add2~13 .shared_arith = "off";

dffeas \adder[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[14]~q ),
	.prn(vcc));
defparam \adder[14] .is_wysiwyg = "true";
defparam \adder[14] .power_up = "low";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\adder[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h00000000000000FF;
defparam \Add2~9 .shared_arith = "off";

dffeas \adder[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Add2~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always15~3_combout ),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\adder[15]~q ),
	.prn(vcc));
defparam \adder[15] .is_wysiwyg = "true";
defparam \adder[15] .power_up = "low";

cyclonev_lcell_comb \always15~0 (
	.dataa(!\adder[15]~q ),
	.datab(!\adder[14]~q ),
	.datac(!\adder[12]~q ),
	.datad(!\adder[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~0 .extended_lut = "off";
defparam \always15~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \always15~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!\adder[10]~q ),
	.datab(!\adder[8]~q ),
	.datac(!\adder[7]~q ),
	.datad(!\adder[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~1 (
	.dataa(!\adder[9]~q ),
	.datab(!\adder[11]~q ),
	.datac(!\always15~0_combout ),
	.datad(!\LessThan3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~1 .extended_lut = "off";
defparam \LessThan3~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \LessThan3~1 .shared_arith = "off";

dffeas inf_64(
	.clk(mac_rx_clock_connection_clk),
	.d(\LessThan3~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\inf_64~q ),
	.prn(vcc));
defparam inf_64.is_wysiwyg = "true";
defparam inf_64.power_up = "low";

cyclonev_lcell_comb \always15~4 (
	.dataa(!\adder[15]~q ),
	.datab(!\adder[14]~q ),
	.datac(!\adder[12]~q ),
	.datad(!\adder[13]~q ),
	.datae(!\cnt_inc~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~4 .extended_lut = "off";
defparam \always15~4 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \always15~4 .shared_arith = "off";

dffeas \frm_max_eq[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always15~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_max_eq[3]~q ),
	.prn(vcc));
defparam \frm_max_eq[3] .is_wysiwyg = "true";
defparam \frm_max_eq[3] .power_up = "low";

cyclonev_lcell_comb \Equal14~0 (
	.dataa(!\adder[10]~q ),
	.datab(!\adder[8]~q ),
	.datac(!\adder[9]~q ),
	.datad(!\adder[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal14~0 .extended_lut = "off";
defparam \Equal14~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \Equal14~0 .shared_arith = "off";

dffeas \frm_max_eq[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal14~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_max_eq[2]~q ),
	.prn(vcc));
defparam \frm_max_eq[2] .is_wysiwyg = "true";
defparam \frm_max_eq[2] .power_up = "low";

cyclonev_lcell_comb \Equal13~0 (
	.dataa(!\adder[7]~q ),
	.datab(!\adder[6]~q ),
	.datac(!\adder[4]~q ),
	.datad(!\adder[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal13~0 .extended_lut = "off";
defparam \Equal13~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \Equal13~0 .shared_arith = "off";

dffeas \frm_max_eq[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal13~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_max_eq[1]~q ),
	.prn(vcc));
defparam \frm_max_eq[1] .is_wysiwyg = "true";
defparam \frm_max_eq[1] .power_up = "low";

cyclonev_lcell_comb \Equal12~0 (
	.dataa(!\adder[0]~q ),
	.datab(!\adder[1]~q ),
	.datac(!\adder[2]~q ),
	.datad(!\adder[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal12~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal12~0 .extended_lut = "off";
defparam \Equal12~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Equal12~0 .shared_arith = "off";

dffeas \frm_max_eq[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal12~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_max_eq[0]~q ),
	.prn(vcc));
defparam \frm_max_eq[0] .is_wysiwyg = "true";
defparam \frm_max_eq[0] .power_up = "low";

cyclonev_lcell_comb \Equal16~0 (
	.dataa(!\frm_max_eq[3]~q ),
	.datab(!\frm_max_eq[2]~q ),
	.datac(!\frm_max_eq[1]~q ),
	.datad(!\frm_max_eq[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal16~0 .extended_lut = "off";
defparam \Equal16~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal16~0 .shared_arith = "off";

dffeas sup_frm_maxv(
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal16~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\sup_frm_maxv~q ),
	.prn(vcc));
defparam sup_frm_maxv.is_wysiwyg = "true";
defparam sup_frm_maxv.power_up = "low";

cyclonev_lcell_comb \always15~2 (
	.dataa(!\inf_64~q ),
	.datab(!\crc_vld[2]~q ),
	.datac(!\sup_frm_maxv~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always15~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always15~2 .extended_lut = "off";
defparam \always15~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always15~2 .shared_arith = "off";

dffeas \frm_lgth_err_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always15~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_lgth_err_reg[0]~q ),
	.prn(vcc));
defparam \frm_lgth_err_reg[0] .is_wysiwyg = "true";
defparam \frm_lgth_err_reg[0] .power_up = "low";

dffeas \frm_lgth_err_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_lgth_err_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_lgth_err_reg[1]~q ),
	.prn(vcc));
defparam \frm_lgth_err_reg[1] .is_wysiwyg = "true";
defparam \frm_lgth_err_reg[1] .power_up = "low";

cyclonev_lcell_comb \end_wr_fifo~0 (
	.dataa(!afull_flag),
	.datab(!\cnt_end_64_user_reg[14]~q ),
	.datac(!\frm_lgth_err_reg[1]~q ),
	.datad(!\rx_en_s[20]~q ),
	.datae(!\rx_en_s[19]~q ),
	.dataf(!\U_SYNC_11|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\end_wr_fifo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \end_wr_fifo~0 .extended_lut = "off";
defparam \end_wr_fifo~0 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \end_wr_fifo~0 .shared_arith = "off";

cyclonev_lcell_comb \end_wr_fifo~1 (
	.dataa(!\fifo_wr~q ),
	.datab(!\U_SYNC_11|std_sync_no_cut|dreg[1]~q ),
	.datac(!\rx_en_s[24]~q ),
	.datad(!\rx_en_s[23]~q ),
	.datae(!\end_wr_fifo~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\end_wr_fifo~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \end_wr_fifo~1 .extended_lut = "off";
defparam \end_wr_fifo~1 .lut_mask = 64'hFFFFFF7FFFFFFF7F;
defparam \end_wr_fifo~1 .shared_arith = "off";

dffeas end_wr_fifo(
	.clk(mac_rx_clock_connection_clk),
	.d(\end_wr_fifo~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\end_wr_fifo~q ),
	.prn(vcc));
defparam end_wr_fifo.is_wysiwyg = "true";
defparam end_wr_fifo.power_up = "low";

cyclonev_lcell_comb \ok_sfd_discard~0 (
	.dataa(!afull_flag),
	.datab(!\no_align_err~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ok_sfd_discard~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ok_sfd_discard~0 .extended_lut = "off";
defparam \ok_sfd_discard~0 .lut_mask = 64'h7777777777777777;
defparam \ok_sfd_discard~0 .shared_arith = "off";

dffeas ok_sfd_discard(
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard~q ),
	.prn(vcc));
defparam ok_sfd_discard.is_wysiwyg = "true";
defparam ok_sfd_discard.power_up = "low";

dffeas \ok_sfd_discard_p[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[0]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[0] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[0] .power_up = "low";

dffeas \ok_sfd_discard_p[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[1]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[1] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[1] .power_up = "low";

dffeas \ok_sfd_discard_p[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[2]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[2] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[2] .power_up = "low";

dffeas \ok_sfd_discard_p[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[3]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[3] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[3] .power_up = "low";

dffeas \ok_sfd_discard_p[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[4]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[4] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[4] .power_up = "low";

dffeas \ok_sfd_discard_p[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[5]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[5] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[5] .power_up = "low";

dffeas \ok_sfd_discard_p[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[6]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[6] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[6] .power_up = "low";

dffeas \ok_sfd_discard_p[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[7]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[7] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[7] .power_up = "low";

dffeas \ok_sfd_discard_p[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[8]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[8] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[8] .power_up = "low";

dffeas \ok_sfd_discard_p[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[9]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[9] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[9] .power_up = "low";

dffeas \ok_sfd_discard_p[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[10]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[10] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[10] .power_up = "low";

dffeas \ok_sfd_discard_p[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[11]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[11] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[11] .power_up = "low";

dffeas \ok_sfd_discard_p[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[12]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[12] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[12] .power_up = "low";

dffeas \ok_sfd_discard_p[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[13]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[13] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[13] .power_up = "low";

dffeas \ok_sfd_discard_p[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[14]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[14] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[14] .power_up = "low";

dffeas \ok_sfd_discard_p[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[14]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[15]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[15] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[15] .power_up = "low";

dffeas \ok_sfd_discard_p[16] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[15]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[16]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[16] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[16] .power_up = "low";

dffeas \ok_sfd_discard_p[17] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[16]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[17]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[17] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[17] .power_up = "low";

dffeas \ok_sfd_discard_p[18] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[17]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[18]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[18] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[18] .power_up = "low";

dffeas \ok_sfd_discard_p[19] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[18]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[19]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[19] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[19] .power_up = "low";

dffeas \ok_sfd_discard_p[20] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[19]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[20]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[20] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[20] .power_up = "low";

dffeas \ok_sfd_discard_p[21] (
	.clk(mac_rx_clock_connection_clk),
	.d(\ok_sfd_discard_p[20]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\ok_sfd_discard_p[21]~q ),
	.prn(vcc));
defparam \ok_sfd_discard_p[21] .is_wysiwyg = "true";
defparam \ok_sfd_discard_p[21] .power_up = "low";

cyclonev_lcell_comb \always14~0 (
	.dataa(!\dest_add_ok[12]~q ),
	.datab(!\user_frm~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~0 .extended_lut = "off";
defparam \always14~0 .lut_mask = 64'h7777777777777777;
defparam \always14~0 .shared_arith = "off";

dffeas frm_to_write(
	.clk(mac_rx_clock_connection_clk),
	.d(\always14~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_to_write~q ),
	.prn(vcc));
defparam frm_to_write.is_wysiwyg = "true";
defparam frm_to_write.power_up = "low";

cyclonev_lcell_comb \always20~3 (
	.dataa(!afull_flag),
	.datab(!\end_wr_fifo~q ),
	.datac(!\ok_sfd_discard_p[21]~q ),
	.datad(!\frm_to_write~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~3 .extended_lut = "off";
defparam \always20~3 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \always20~3 .shared_arith = "off";

dffeas start_wr_fifo(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\start_wr_fifo~q ),
	.prn(vcc));
defparam start_wr_fifo.is_wysiwyg = "true";
defparam start_wr_fifo.power_up = "low";

cyclonev_lcell_comb \always20~4 (
	.dataa(!\start_wr_fifo~q ),
	.datab(!\fifo_wr_wait~q ),
	.datac(!\fifo_wr~q ),
	.datad(!\end_wr_fifo~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~4 .extended_lut = "off";
defparam \always20~4 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \always20~4 .shared_arith = "off";

dffeas fifo_wr_wait(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\fifo_wr_wait~q ),
	.prn(vcc));
defparam fifo_wr_wait.is_wysiwyg = "true";
defparam fifo_wr_wait.power_up = "low";

cyclonev_lcell_comb \always20~5 (
	.dataa(!\start_wr_fifo~q ),
	.datab(!\fifo_wr_wait~q ),
	.datac(!\fifo_wr~q ),
	.datad(!\end_wr_fifo~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~5 .extended_lut = "off";
defparam \always20~5 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \always20~5 .shared_arith = "off";

dffeas fifo_wr(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclonev_lcell_comb \user_p_lgth_inf_46_reg~2 (
	.dataa(!\crc_vld[5]~q ),
	.datab(!\user_p_lgth_inf_46_reg[1]~q ),
	.datac(!\user_p_lgth_inf_46_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_p_lgth_inf_46_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_p_lgth_inf_46_reg~2 .extended_lut = "off";
defparam \user_p_lgth_inf_46_reg~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \user_p_lgth_inf_46_reg~2 .shared_arith = "off";

dffeas \user_p_lgth_inf_46_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\user_p_lgth_inf_46_reg~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\user_p_lgth_inf_46_reg[1]~q ),
	.prn(vcc));
defparam \user_p_lgth_inf_46_reg[1] .is_wysiwyg = "true";
defparam \user_p_lgth_inf_46_reg[1] .power_up = "low";

cyclonev_lcell_comb \always20~8 (
	.dataa(!\fifo_wr~q ),
	.datab(!\end_wr_fifo~q ),
	.datac(!\stat_wr_wait~q ),
	.datad(!\user_p_lgth_inf_46_reg[1]~q ),
	.datae(!\U_CRC|eof_dly[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~8 .extended_lut = "off";
defparam \always20~8 .lut_mask = 64'hF377FFFFF377FFFF;
defparam \always20~8 .shared_arith = "off";

dffeas stat_wr(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\stat_wr~q ),
	.prn(vcc));
defparam stat_wr.is_wysiwyg = "true";
defparam stat_wr.power_up = "low";

cyclonev_lcell_comb \always20~7 (
	.dataa(!\fifo_wr~q ),
	.datab(!\end_wr_fifo~q ),
	.datac(!\stat_wr_wait~q ),
	.datad(!\stat_wr~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~7 .extended_lut = "off";
defparam \always20~7 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \always20~7 .shared_arith = "off";

dffeas stat_wr_wait(
	.clk(mac_rx_clock_connection_clk),
	.d(\always20~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\stat_wr_wait~q ),
	.prn(vcc));
defparam stat_wr_wait.is_wysiwyg = "true";
defparam stat_wr_wait.power_up = "low";

cyclonev_lcell_comb \rx_stat_wren_s~0 (
	.dataa(!\fifo_wr~q ),
	.datab(!\end_wr_fifo~q ),
	.datac(!\rx_stat_wren_s[0]~q ),
	.datad(!\stat_wr_wait~q ),
	.datae(!\user_p_lgth_inf_46_reg[1]~q ),
	.dataf(!\U_CRC|eof_dly[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_wren_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_wren_s~0 .extended_lut = "off";
defparam \rx_stat_wren_s~0 .lut_mask = 64'hFF3F7F7FFFFFFFFF;
defparam \rx_stat_wren_s~0 .shared_arith = "off";

dffeas \rx_stat_wren_s[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[0]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[0] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[0] .power_up = "low";

dffeas \rx_stat_wren_s[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[1]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[1] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[1] .power_up = "low";

dffeas \rx_stat_wren_s[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[2]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[2] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[2] .power_up = "low";

dffeas \rx_stat_wren_s[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[3]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[3] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[3] .power_up = "low";

dffeas \rx_stat_wren_s[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[4]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[4] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[4] .power_up = "low";

dffeas \rx_stat_wren_s[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[5]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[5] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[5] .power_up = "low";

dffeas \rx_stat_wren_s[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[6]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[6] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[6] .power_up = "low";

dffeas \rx_stat_wren_s[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[7]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[7] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[7] .power_up = "low";

dffeas \rx_stat_wren_s[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[8]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[8] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[8] .power_up = "low";

dffeas \rx_stat_wren_s[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[9]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[9] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[9] .power_up = "low";

dffeas \rx_stat_wren_s[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[10]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[10] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[10] .power_up = "low";

dffeas \rx_stat_wren_s[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_stat_wren_s[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_stat_wren_s[11]~q ),
	.prn(vcc));
defparam \rx_stat_wren_s[11] .is_wysiwyg = "true";
defparam \rx_stat_wren_s[11] .power_up = "low";

cyclonev_lcell_comb \current_frame~0 (
	.dataa(!\current_frame~q ),
	.datab(!\start_wr_fifo~q ),
	.datac(!\rx_stat_wren_s[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_frame~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_frame~0 .extended_lut = "off";
defparam \current_frame~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \current_frame~0 .shared_arith = "off";

dffeas current_frame(
	.clk(mac_rx_clock_connection_clk),
	.d(\current_frame~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_frame~q ),
	.prn(vcc));
defparam current_frame.is_wysiwyg = "true";
defparam current_frame.power_up = "low";

cyclonev_lcell_comb \sleep_mode_ena~0 (
	.dataa(!\sleep_mode_ena~q ),
	.datab(!\current_frame~q ),
	.datac(!\U_SYNC_3|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sleep_mode_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sleep_mode_ena~0 .extended_lut = "off";
defparam \sleep_mode_ena~0 .lut_mask = 64'h4747474747474747;
defparam \sleep_mode_ena~0 .shared_arith = "off";

dffeas sleep_mode_ena(
	.clk(mac_rx_clock_connection_clk),
	.d(\sleep_mode_ena~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sleep_mode_ena~q ),
	.prn(vcc));
defparam sleep_mode_ena.is_wysiwyg = "true";
defparam sleep_mode_ena.power_up = "low";

cyclonev_lcell_comb \rx_stat_wren~0 (
	.dataa(!\rx_stat_wren_s[9]~q ),
	.datab(!rxclk_ena),
	.datac(!\sleep_mode_ena~q ),
	.datad(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_wren~0 .extended_lut = "off";
defparam \rx_stat_wren~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \rx_stat_wren~0 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[0]~1 (
	.dataa(!\user_length[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[0]~1 .extended_lut = "off";
defparam \payload_length[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[0]~0 (
	.dataa(!rxclk_ena),
	.datab(!\rx_en_s[12]~q ),
	.datac(!\rx_en_s[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[0]~0 .extended_lut = "off";
defparam \payload_length[0]~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \payload_length[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[1]~2 (
	.dataa(!\user_length[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[1]~2 .extended_lut = "off";
defparam \payload_length[1]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[2]~3 (
	.dataa(!\user_length[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[2]~3 .extended_lut = "off";
defparam \payload_length[2]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[3]~4 (
	.dataa(!\user_length[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[3]~4 .extended_lut = "off";
defparam \payload_length[3]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[4]~5 (
	.dataa(!\user_length[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[4]~5 .extended_lut = "off";
defparam \payload_length[4]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[5]~6 (
	.dataa(!\user_length[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[5]~6 .extended_lut = "off";
defparam \payload_length[5]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[6]~7 (
	.dataa(!\user_length[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[6]~7 .extended_lut = "off";
defparam \payload_length[6]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[7]~8 (
	.dataa(!\user_length[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[7]~8 .extended_lut = "off";
defparam \payload_length[7]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[8]~9 (
	.dataa(!\user_length[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[8]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[8]~9 .extended_lut = "off";
defparam \payload_length[8]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[8]~9 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[9]~10 (
	.dataa(!\user_length[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[9]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[9]~10 .extended_lut = "off";
defparam \payload_length[9]~10 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[9]~10 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[10]~11 (
	.dataa(!\user_length[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[10]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[10]~11 .extended_lut = "off";
defparam \payload_length[10]~11 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[10]~11 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[11]~12 (
	.dataa(!\user_length[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[11]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[11]~12 .extended_lut = "off";
defparam \payload_length[11]~12 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[11]~12 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[12]~13 (
	.dataa(!\user_length[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[12]~13 .extended_lut = "off";
defparam \payload_length[12]~13 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[12]~13 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[13]~14 (
	.dataa(!\user_length[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[13]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[13]~14 .extended_lut = "off";
defparam \payload_length[13]~14 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[13]~14 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[14]~15 (
	.dataa(!\user_length[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[14]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[14]~15 .extended_lut = "off";
defparam \payload_length[14]~15 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[14]~15 .shared_arith = "off";

cyclonev_lcell_comb \payload_length[15]~16 (
	.dataa(!\user_length[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\payload_length[15]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \payload_length[15]~16 .extended_lut = "off";
defparam \payload_length[15]~16 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \payload_length[15]~16 .shared_arith = "off";

cyclonev_lcell_comb \always20~0 (
	.dataa(!rxclk_ena),
	.datab(!\sleep_mode_ena~q ),
	.datac(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datad(!\start_wr_fifo~q ),
	.datae(!\fifo_wr_wait~q ),
	.dataf(!\fifo_wr~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~0 .extended_lut = "off";
defparam \always20~0 .lut_mask = 64'hFFFFFDFFFFFFFFFF;
defparam \always20~0 .shared_arith = "off";

cyclonev_lcell_comb \always20~1 (
	.dataa(!\fifo_wr~q ),
	.datab(!\end_wr_fifo~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~1 .extended_lut = "off";
defparam \always20~1 .lut_mask = 64'h7777777777777777;
defparam \always20~1 .shared_arith = "off";

dffeas \gm_rx_col_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SYNC_13|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\gm_rx_col_reg[0]~q ),
	.prn(vcc));
defparam \gm_rx_col_reg[0] .is_wysiwyg = "true";
defparam \gm_rx_col_reg[0] .power_up = "low";

dffeas \gm_rx_col_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\gm_rx_col_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\gm_rx_col_reg[1]~q ),
	.prn(vcc));
defparam \gm_rx_col_reg[1] .is_wysiwyg = "true";
defparam \gm_rx_col_reg[1] .power_up = "low";

dffeas \gm_rx_col_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\gm_rx_col_reg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\gm_rx_col_reg[2]~q ),
	.prn(vcc));
defparam \gm_rx_col_reg[2] .is_wysiwyg = "true";
defparam \gm_rx_col_reg[2] .power_up = "low";

dffeas \gm_rx_col_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\gm_rx_col_reg[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\gm_rx_col_reg[3]~q ),
	.prn(vcc));
defparam \gm_rx_col_reg[3] .is_wysiwyg = "true";
defparam \gm_rx_col_reg[3] .power_up = "low";

cyclonev_lcell_comb \col_int~0 (
	.dataa(!en),
	.datab(!\col_int~q ),
	.datac(!\U_SYNC_1|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_10|std_sync_no_cut|dreg[1]~q ),
	.datae(!\gm_rx_col_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\col_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_int~0 .extended_lut = "off";
defparam \col_int~0 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \col_int~0 .shared_arith = "off";

dffeas col_int(
	.clk(mac_rx_clock_connection_clk),
	.d(\col_int~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\col_int~q ),
	.prn(vcc));
defparam col_int.is_wysiwyg = "true";
defparam col_int.power_up = "low";

dffeas \col_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_int~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[0]~q ),
	.prn(vcc));
defparam \col_reg[0] .is_wysiwyg = "true";
defparam \col_reg[0] .power_up = "low";

dffeas \col_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[1]~q ),
	.prn(vcc));
defparam \col_reg[1] .is_wysiwyg = "true";
defparam \col_reg[1] .power_up = "low";

dffeas \col_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[2]~q ),
	.prn(vcc));
defparam \col_reg[2] .is_wysiwyg = "true";
defparam \col_reg[2] .power_up = "low";

dffeas \col_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[3]~q ),
	.prn(vcc));
defparam \col_reg[3] .is_wysiwyg = "true";
defparam \col_reg[3] .power_up = "low";

dffeas \col_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[4]~q ),
	.prn(vcc));
defparam \col_reg[4] .is_wysiwyg = "true";
defparam \col_reg[4] .power_up = "low";

dffeas \col_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[5]~q ),
	.prn(vcc));
defparam \col_reg[5] .is_wysiwyg = "true";
defparam \col_reg[5] .power_up = "low";

dffeas \col_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[6]~q ),
	.prn(vcc));
defparam \col_reg[6] .is_wysiwyg = "true";
defparam \col_reg[6] .power_up = "low";

dffeas \col_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[7]~q ),
	.prn(vcc));
defparam \col_reg[7] .is_wysiwyg = "true";
defparam \col_reg[7] .power_up = "low";

dffeas \col_reg[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[8]~q ),
	.prn(vcc));
defparam \col_reg[8] .is_wysiwyg = "true";
defparam \col_reg[8] .power_up = "low";

dffeas \col_reg[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[9]~q ),
	.prn(vcc));
defparam \col_reg[9] .is_wysiwyg = "true";
defparam \col_reg[9] .power_up = "low";

dffeas \col_reg[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[10]~q ),
	.prn(vcc));
defparam \col_reg[10] .is_wysiwyg = "true";
defparam \col_reg[10] .power_up = "low";

dffeas \col_reg[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[11]~q ),
	.prn(vcc));
defparam \col_reg[11] .is_wysiwyg = "true";
defparam \col_reg[11] .power_up = "low";

dffeas \col_reg[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[12]~q ),
	.prn(vcc));
defparam \col_reg[12] .is_wysiwyg = "true";
defparam \col_reg[12] .power_up = "low";

dffeas \col_reg[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[13]~q ),
	.prn(vcc));
defparam \col_reg[13] .is_wysiwyg = "true";
defparam \col_reg[13] .power_up = "low";

dffeas \col_reg[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[14]~q ),
	.prn(vcc));
defparam \col_reg[14] .is_wysiwyg = "true";
defparam \col_reg[14] .power_up = "low";

dffeas \col_reg[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[14]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[15]~q ),
	.prn(vcc));
defparam \col_reg[15] .is_wysiwyg = "true";
defparam \col_reg[15] .power_up = "low";

dffeas \col_reg[16] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[15]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[16]~q ),
	.prn(vcc));
defparam \col_reg[16] .is_wysiwyg = "true";
defparam \col_reg[16] .power_up = "low";

dffeas \col_reg[17] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[16]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[17]~q ),
	.prn(vcc));
defparam \col_reg[17] .is_wysiwyg = "true";
defparam \col_reg[17] .power_up = "low";

dffeas \col_reg[18] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[17]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[18]~q ),
	.prn(vcc));
defparam \col_reg[18] .is_wysiwyg = "true";
defparam \col_reg[18] .power_up = "low";

dffeas \col_reg[19] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[18]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[19]~q ),
	.prn(vcc));
defparam \col_reg[19] .is_wysiwyg = "true";
defparam \col_reg[19] .power_up = "low";

dffeas \col_reg[20] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[19]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[20]~q ),
	.prn(vcc));
defparam \col_reg[20] .is_wysiwyg = "true";
defparam \col_reg[20] .power_up = "low";

dffeas \col_reg[21] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[20]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[21]~q ),
	.prn(vcc));
defparam \col_reg[21] .is_wysiwyg = "true";
defparam \col_reg[21] .power_up = "low";

dffeas \col_reg[22] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[21]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[22]~q ),
	.prn(vcc));
defparam \col_reg[22] .is_wysiwyg = "true";
defparam \col_reg[22] .power_up = "low";

dffeas \col_reg[23] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[22]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[23]~q ),
	.prn(vcc));
defparam \col_reg[23] .is_wysiwyg = "true";
defparam \col_reg[23] .power_up = "low";

dffeas \col_reg[24] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[23]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[24]~q ),
	.prn(vcc));
defparam \col_reg[24] .is_wysiwyg = "true";
defparam \col_reg[24] .power_up = "low";

dffeas \col_reg[25] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[24]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[25]~q ),
	.prn(vcc));
defparam \col_reg[25] .is_wysiwyg = "true";
defparam \col_reg[25] .power_up = "low";

dffeas \col_reg[26] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[25]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[26]~q ),
	.prn(vcc));
defparam \col_reg[26] .is_wysiwyg = "true";
defparam \col_reg[26] .power_up = "low";

dffeas \col_reg[27] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[26]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[27]~q ),
	.prn(vcc));
defparam \col_reg[27] .is_wysiwyg = "true";
defparam \col_reg[27] .power_up = "low";

dffeas \col_reg[28] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[27]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[28]~q ),
	.prn(vcc));
defparam \col_reg[28] .is_wysiwyg = "true";
defparam \col_reg[28] .power_up = "low";

dffeas \col_reg[29] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[28]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[29]~q ),
	.prn(vcc));
defparam \col_reg[29] .is_wysiwyg = "true";
defparam \col_reg[29] .power_up = "low";

dffeas \col_reg[30] (
	.clk(mac_rx_clock_connection_clk),
	.d(\col_reg[29]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\col_reg[30]~q ),
	.prn(vcc));
defparam \col_reg[30] .is_wysiwyg = "true";
defparam \col_reg[30] .power_up = "low";

cyclonev_lcell_comb \rx_stat_data_s~0 (
	.dataa(!rx_stat_data_s_5),
	.datab(!\rx_stat_wren_s[2]~q ),
	.datac(!\col_reg[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_data_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_data_s~0 .extended_lut = "off";
defparam \rx_stat_data_s~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \rx_stat_data_s~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~0 (
	.dataa(!\user_length[8]~q ),
	.datab(!\user_length[9]~q ),
	.datac(!\user_length[10]~q ),
	.datad(!\adder[10]~q ),
	.datae(!\adder[8]~q ),
	.dataf(!\adder[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~0 .extended_lut = "off";
defparam \Equal17~0 .lut_mask = 64'h6996966996696996;
defparam \Equal17~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~1 (
	.dataa(!\user_length[5]~q ),
	.datab(!\user_length[6]~q ),
	.datac(!\user_length[7]~q ),
	.datad(!\adder[7]~q ),
	.datae(!\adder[6]~q ),
	.dataf(!\adder[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~1 .extended_lut = "off";
defparam \Equal17~1 .lut_mask = 64'h6996966996696996;
defparam \Equal17~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~2 (
	.dataa(!\user_length[0]~q ),
	.datab(!\user_length[1]~q ),
	.datac(!\adder[11]~q ),
	.datad(!\adder[0]~q ),
	.datae(!\adder[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~2 .extended_lut = "off";
defparam \Equal17~2 .lut_mask = 64'hF6F9F9F6F6F9F9F6;
defparam \Equal17~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~3 (
	.dataa(!\user_length[2]~q ),
	.datab(!\user_length[3]~q ),
	.datac(!\user_length[4]~q ),
	.datad(!\adder[2]~q ),
	.datae(!\adder[3]~q ),
	.dataf(!\adder[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~3 .extended_lut = "off";
defparam \Equal17~3 .lut_mask = 64'h6996966996696996;
defparam \Equal17~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal17~4 (
	.dataa(!\always15~0_combout ),
	.datab(!\Equal17~0_combout ),
	.datac(!\Equal17~1_combout ),
	.datad(!\Equal17~2_combout ),
	.datae(!\Equal17~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal17~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal17~4 .extended_lut = "off";
defparam \Equal17~4 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \Equal17~4 .shared_arith = "off";

cyclonev_lcell_comb \frm_length_error~0 (
	.dataa(!\user_length[9]~q ),
	.datab(!\user_length[10]~q ),
	.datac(!\rx_en_s[9]~q ),
	.datad(!\rx_en_s[8]~q ),
	.datae(!\always15~1_combout ),
	.dataf(!\user_p_lgth_inf_46_reg~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_length_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_length_error~0 .extended_lut = "off";
defparam \frm_length_error~0 .lut_mask = 64'hFF7FFFFFDF5FFFFF;
defparam \frm_length_error~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_length_error~1 (
	.dataa(!\end_wr_fifo~q ),
	.datab(!\rx_en_s[9]~q ),
	.datac(!\frm_length_error~q ),
	.datad(!\rx_en_s[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_length_error~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_length_error~1 .extended_lut = "off";
defparam \frm_length_error~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \frm_length_error~1 .shared_arith = "off";

cyclonev_lcell_comb \frm_length_error~2 (
	.dataa(!\U_SYNC_7|std_sync_no_cut|dreg[1]~q ),
	.datab(!\Equal17~4_combout ),
	.datac(!\user_p_lgth_inf_46_reg~0_combout ),
	.datad(!\frm_length_error~0_combout ),
	.datae(!\frm_length_error~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_length_error~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_length_error~2 .extended_lut = "off";
defparam \frm_length_error~2 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \frm_length_error~2 .shared_arith = "off";

dffeas frm_length_error(
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_length_error~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_length_error~q ),
	.prn(vcc));
defparam frm_length_error.is_wysiwyg = "true";
defparam frm_length_error.power_up = "low";

cyclonev_lcell_comb \frm_lgth_err_s_reg~0 (
	.dataa(!\frm_lgth_err_s_reg~q ),
	.datab(!\inf_64~q ),
	.datac(!\crc_vld[2]~q ),
	.datad(!\sup_frm_maxv~q ),
	.datae(!\frm_length_error~q ),
	.dataf(!\crc_vld[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_lgth_err_s_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_lgth_err_s_reg~0 .extended_lut = "off";
defparam \frm_lgth_err_s_reg~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \frm_lgth_err_s_reg~0 .shared_arith = "off";

dffeas frm_lgth_err_s_reg(
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_lgth_err_s_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_lgth_err_s_reg~q ),
	.prn(vcc));
defparam frm_lgth_err_s_reg.is_wysiwyg = "true";
defparam frm_lgth_err_s_reg.power_up = "low";

cyclonev_lcell_comb \rx_stat_data_s~1 (
	.dataa(!rx_stat_data_s_0),
	.datab(!\rx_stat_wren_s[2]~q ),
	.datac(!\frm_lgth_err_s_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_data_s~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_data_s~1 .extended_lut = "off";
defparam \rx_stat_data_s~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \rx_stat_data_s~1 .shared_arith = "off";

dffeas \crc_ok[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_CRC|crc_ok~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_ok[1]~q ),
	.prn(vcc));
defparam \crc_ok[1] .is_wysiwyg = "true";
defparam \crc_ok[1] .power_up = "low";

dffeas \crc_ok[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_ok[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_ok[2]~q ),
	.prn(vcc));
defparam \crc_ok[2] .is_wysiwyg = "true";
defparam \crc_ok[2] .power_up = "low";

dffeas \crc_ok[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_ok[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_ok[3]~q ),
	.prn(vcc));
defparam \crc_ok[3] .is_wysiwyg = "true";
defparam \crc_ok[3] .power_up = "low";

dffeas \crc_ok[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\crc_ok[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\crc_ok[4]~q ),
	.prn(vcc));
defparam \crc_ok[4] .is_wysiwyg = "true";
defparam \crc_ok[4] .power_up = "low";

cyclonev_lcell_comb \rx_stat_data_s~2 (
	.dataa(!rx_stat_data_s_1),
	.datab(!\rx_stat_wren_s[2]~q ),
	.datac(!\crc_vld[4]~q ),
	.datad(!\crc_ok[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_data_s~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_data_s~2 .extended_lut = "off";
defparam \rx_stat_data_s~2 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \rx_stat_data_s~2 .shared_arith = "off";

cyclonev_lcell_comb \rx_a_full_s~0 (
	.dataa(!afull_flag),
	.datab(!\rx_stat_wren_s[9]~q ),
	.datac(!\start_wr_fifo~q ),
	.datad(!\fifo_wr_wait~q ),
	.datae(!\fifo_wr~q ),
	.dataf(!\rx_a_full_s~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_a_full_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_a_full_s~0 .extended_lut = "off";
defparam \rx_a_full_s~0 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \rx_a_full_s~0 .shared_arith = "off";

dffeas rx_a_full_s(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_a_full_s~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_a_full_s~q ),
	.prn(vcc));
defparam rx_a_full_s.is_wysiwyg = "true";
defparam rx_a_full_s.power_up = "low";

cyclonev_lcell_comb \rx_stat_data_s~3 (
	.dataa(!rx_stat_data_s_2),
	.datab(!\rx_stat_wren_s[2]~q ),
	.datac(!\rx_a_full_s~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_data_s~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_data_s~3 .extended_lut = "off";
defparam \rx_stat_data_s~3 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \rx_stat_data_s~3 .shared_arith = "off";

cyclonev_lcell_comb \rx_err_s~0 (
	.dataa(!\enable_rx_reg3~q ),
	.datab(!en),
	.datac(!err),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_err_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_err_s~0 .extended_lut = "off";
defparam \rx_err_s~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \rx_err_s~0 .shared_arith = "off";

dffeas \rx_err_s[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[0]~q ),
	.prn(vcc));
defparam \rx_err_s[0] .is_wysiwyg = "true";
defparam \rx_err_s[0] .power_up = "low";

dffeas \rx_err_s[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[1]~q ),
	.prn(vcc));
defparam \rx_err_s[1] .is_wysiwyg = "true";
defparam \rx_err_s[1] .power_up = "low";

dffeas \rx_err_s[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[2]~q ),
	.prn(vcc));
defparam \rx_err_s[2] .is_wysiwyg = "true";
defparam \rx_err_s[2] .power_up = "low";

dffeas \rx_err_s[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[3]~q ),
	.prn(vcc));
defparam \rx_err_s[3] .is_wysiwyg = "true";
defparam \rx_err_s[3] .power_up = "low";

dffeas \rx_err_s[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[4]~q ),
	.prn(vcc));
defparam \rx_err_s[4] .is_wysiwyg = "true";
defparam \rx_err_s[4] .power_up = "low";

dffeas \rx_err_s[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[5]~q ),
	.prn(vcc));
defparam \rx_err_s[5] .is_wysiwyg = "true";
defparam \rx_err_s[5] .power_up = "low";

dffeas \rx_err_s[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[6]~q ),
	.prn(vcc));
defparam \rx_err_s[6] .is_wysiwyg = "true";
defparam \rx_err_s[6] .power_up = "low";

dffeas \rx_err_s[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[7]~q ),
	.prn(vcc));
defparam \rx_err_s[7] .is_wysiwyg = "true";
defparam \rx_err_s[7] .power_up = "low";

dffeas \rx_err_s[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[8]~q ),
	.prn(vcc));
defparam \rx_err_s[8] .is_wysiwyg = "true";
defparam \rx_err_s[8] .power_up = "low";

dffeas \rx_err_s[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[9]~q ),
	.prn(vcc));
defparam \rx_err_s[9] .is_wysiwyg = "true";
defparam \rx_err_s[9] .power_up = "low";

dffeas \rx_err_s[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[10]~q ),
	.prn(vcc));
defparam \rx_err_s[10] .is_wysiwyg = "true";
defparam \rx_err_s[10] .power_up = "low";

dffeas \rx_err_s[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[11]~q ),
	.prn(vcc));
defparam \rx_err_s[11] .is_wysiwyg = "true";
defparam \rx_err_s[11] .power_up = "low";

dffeas \rx_err_s[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[12]~q ),
	.prn(vcc));
defparam \rx_err_s[12] .is_wysiwyg = "true";
defparam \rx_err_s[12] .power_up = "low";

dffeas \rx_err_s[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[13]~q ),
	.prn(vcc));
defparam \rx_err_s[13] .is_wysiwyg = "true";
defparam \rx_err_s[13] .power_up = "low";

dffeas \rx_err_s[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[14]~q ),
	.prn(vcc));
defparam \rx_err_s[14] .is_wysiwyg = "true";
defparam \rx_err_s[14] .power_up = "low";

dffeas \rx_err_s[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[14]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[15]~q ),
	.prn(vcc));
defparam \rx_err_s[15] .is_wysiwyg = "true";
defparam \rx_err_s[15] .power_up = "low";

dffeas \rx_err_s[16] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[15]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[16]~q ),
	.prn(vcc));
defparam \rx_err_s[16] .is_wysiwyg = "true";
defparam \rx_err_s[16] .power_up = "low";

dffeas \rx_err_s[17] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[16]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[17]~q ),
	.prn(vcc));
defparam \rx_err_s[17] .is_wysiwyg = "true";
defparam \rx_err_s[17] .power_up = "low";

dffeas \rx_err_s[18] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[17]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[18]~q ),
	.prn(vcc));
defparam \rx_err_s[18] .is_wysiwyg = "true";
defparam \rx_err_s[18] .power_up = "low";

dffeas \rx_err_s[19] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[18]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[19]~q ),
	.prn(vcc));
defparam \rx_err_s[19] .is_wysiwyg = "true";
defparam \rx_err_s[19] .power_up = "low";

dffeas \rx_err_s[20] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[19]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[20]~q ),
	.prn(vcc));
defparam \rx_err_s[20] .is_wysiwyg = "true";
defparam \rx_err_s[20] .power_up = "low";

dffeas \rx_err_s[21] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[20]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[21]~q ),
	.prn(vcc));
defparam \rx_err_s[21] .is_wysiwyg = "true";
defparam \rx_err_s[21] .power_up = "low";

dffeas \rx_err_s[22] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[21]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[22]~q ),
	.prn(vcc));
defparam \rx_err_s[22] .is_wysiwyg = "true";
defparam \rx_err_s[22] .power_up = "low";

dffeas \rx_err_s[23] (
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_s[22]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_s[23]~q ),
	.prn(vcc));
defparam \rx_err_s[23] .is_wysiwyg = "true";
defparam \rx_err_s[23] .power_up = "low";

cyclonev_lcell_comb \rx_err_latched_temp~0 (
	.dataa(!\rx_en_s[24]~q ),
	.datab(!\rx_en_s[25]~q ),
	.datac(!\rx_err_latched_temp~q ),
	.datad(!\rx_err_s[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_err_latched_temp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_err_latched_temp~0 .extended_lut = "off";
defparam \rx_err_latched_temp~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \rx_err_latched_temp~0 .shared_arith = "off";

dffeas rx_err_latched_temp(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_latched_temp~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_latched_temp~q ),
	.prn(vcc));
defparam rx_err_latched_temp.is_wysiwyg = "true";
defparam rx_err_latched_temp.power_up = "low";

dffeas \frm_type_ok_s[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_type_ok_s[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_type_ok_s[1]~q ),
	.prn(vcc));
defparam \frm_type_ok_s[1] .is_wysiwyg = "true";
defparam \frm_type_ok_s[1] .power_up = "low";

cyclonev_lcell_comb \frm_ok~0 (
	.dataa(!\rx_en_s[24]~q ),
	.datab(!\rx_en_s[25]~q ),
	.datac(!\frm_ok~q ),
	.datad(!\frm_type_ok_s[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_ok~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_ok~0 .extended_lut = "off";
defparam \frm_ok~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \frm_ok~0 .shared_arith = "off";

dffeas frm_ok(
	.clk(mac_rx_clock_connection_clk),
	.d(\frm_ok~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\frm_ok~q ),
	.prn(vcc));
defparam frm_ok.is_wysiwyg = "true";
defparam frm_ok.power_up = "low";

cyclonev_lcell_comb \rx_err_latched~0 (
	.dataa(!\rx_err_latched~q ),
	.datab(!\rx_en_s[24]~q ),
	.datac(!\rx_en_s[25]~q ),
	.datad(!\rx_err_latched_temp~q ),
	.datae(!\frm_ok~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_err_latched~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_err_latched~0 .extended_lut = "off";
defparam \rx_err_latched~0 .lut_mask = 64'hF3FF77FFF3FF77FF;
defparam \rx_err_latched~0 .shared_arith = "off";

dffeas rx_err_latched(
	.clk(mac_rx_clock_connection_clk),
	.d(\rx_err_latched~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rx_err_latched~q ),
	.prn(vcc));
defparam rx_err_latched.is_wysiwyg = "true";
defparam rx_err_latched.power_up = "low";

cyclonev_lcell_comb \rx_stat_data_s~4 (
	.dataa(!rx_stat_data_s_3),
	.datab(!\rx_stat_wren_s[2]~q ),
	.datac(!\rx_err_latched~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_stat_data_s~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_stat_data_s~4 .extended_lut = "off";
defparam \rx_stat_data_s~4 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \rx_stat_data_s~4 .shared_arith = "off";

cyclonev_lcell_comb \always20~2 (
	.dataa(!\start_wr_fifo~q ),
	.datab(!\fifo_wr_wait~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~2 .extended_lut = "off";
defparam \always20~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always20~2 .shared_arith = "off";

cyclonev_lcell_comb \always10~15 (
	.dataa(!\rxd_8[0]~q ),
	.datab(!\ok_sfd_p[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~15 .extended_lut = "off";
defparam \always10~15 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always10~15 .shared_arith = "off";

dffeas \unicast_add_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\always10~15_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[0]~q ),
	.prn(vcc));
defparam \unicast_add_reg[0] .is_wysiwyg = "true";
defparam \unicast_add_reg[0] .power_up = "low";

dffeas \unicast_add_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[1]~q ),
	.prn(vcc));
defparam \unicast_add_reg[1] .is_wysiwyg = "true";
defparam \unicast_add_reg[1] .power_up = "low";

dffeas \unicast_add_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[2]~q ),
	.prn(vcc));
defparam \unicast_add_reg[2] .is_wysiwyg = "true";
defparam \unicast_add_reg[2] .power_up = "low";

dffeas \unicast_add_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[3]~q ),
	.prn(vcc));
defparam \unicast_add_reg[3] .is_wysiwyg = "true";
defparam \unicast_add_reg[3] .power_up = "low";

dffeas \unicast_add_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[4]~q ),
	.prn(vcc));
defparam \unicast_add_reg[4] .is_wysiwyg = "true";
defparam \unicast_add_reg[4] .power_up = "low";

dffeas \unicast_add_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[5]~q ),
	.prn(vcc));
defparam \unicast_add_reg[5] .is_wysiwyg = "true";
defparam \unicast_add_reg[5] .power_up = "low";

dffeas \unicast_add_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[6]~q ),
	.prn(vcc));
defparam \unicast_add_reg[6] .is_wysiwyg = "true";
defparam \unicast_add_reg[6] .power_up = "low";

dffeas \unicast_add_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[7]~q ),
	.prn(vcc));
defparam \unicast_add_reg[7] .is_wysiwyg = "true";
defparam \unicast_add_reg[7] .power_up = "low";

dffeas \unicast_add_reg[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[8]~q ),
	.prn(vcc));
defparam \unicast_add_reg[8] .is_wysiwyg = "true";
defparam \unicast_add_reg[8] .power_up = "low";

dffeas \unicast_add_reg[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[9]~q ),
	.prn(vcc));
defparam \unicast_add_reg[9] .is_wysiwyg = "true";
defparam \unicast_add_reg[9] .power_up = "low";

dffeas \unicast_add_reg[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[10]~q ),
	.prn(vcc));
defparam \unicast_add_reg[10] .is_wysiwyg = "true";
defparam \unicast_add_reg[10] .power_up = "low";

dffeas \unicast_add_reg[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[11]~q ),
	.prn(vcc));
defparam \unicast_add_reg[11] .is_wysiwyg = "true";
defparam \unicast_add_reg[11] .power_up = "low";

dffeas \unicast_add_reg[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[12]~q ),
	.prn(vcc));
defparam \unicast_add_reg[12] .is_wysiwyg = "true";
defparam \unicast_add_reg[12] .power_up = "low";

dffeas \unicast_add_reg[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[13]~q ),
	.prn(vcc));
defparam \unicast_add_reg[13] .is_wysiwyg = "true";
defparam \unicast_add_reg[13] .power_up = "low";

dffeas \unicast_add_reg[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[14]~q ),
	.prn(vcc));
defparam \unicast_add_reg[14] .is_wysiwyg = "true";
defparam \unicast_add_reg[14] .power_up = "low";

dffeas \unicast_add_reg[15] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[14]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[15]~q ),
	.prn(vcc));
defparam \unicast_add_reg[15] .is_wysiwyg = "true";
defparam \unicast_add_reg[15] .power_up = "low";

dffeas \unicast_add_reg[16] (
	.clk(mac_rx_clock_connection_clk),
	.d(\unicast_add_reg[15]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\unicast_add_reg[16]~q ),
	.prn(vcc));
defparam \unicast_add_reg[16] .is_wysiwyg = "true";
defparam \unicast_add_reg[16] .power_up = "low";

cyclonev_lcell_comb \broad_add_reg~0 (
	.dataa(!\always20~2_combout ),
	.datab(!\broad_add_reg~q ),
	.datac(!\broad_sub[0]~q ),
	.datad(!\ok_sfd_p[6]~q ),
	.datae(!\always9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\broad_add_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \broad_add_reg~0 .extended_lut = "off";
defparam \broad_add_reg~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \broad_add_reg~0 .shared_arith = "off";

dffeas broad_add_reg(
	.clk(mac_rx_clock_connection_clk),
	.d(\broad_add_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\broad_add_reg~q ),
	.prn(vcc));
defparam broad_add_reg.is_wysiwyg = "true";
defparam broad_add_reg.power_up = "low";

dffeas \multicast_add_reg[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_en[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[0]~q ),
	.prn(vcc));
defparam \multicast_add_reg[0] .is_wysiwyg = "true";
defparam \multicast_add_reg[0] .power_up = "low";

dffeas \multicast_add_reg[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[1]~q ),
	.prn(vcc));
defparam \multicast_add_reg[1] .is_wysiwyg = "true";
defparam \multicast_add_reg[1] .power_up = "low";

dffeas \multicast_add_reg[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[2]~q ),
	.prn(vcc));
defparam \multicast_add_reg[2] .is_wysiwyg = "true";
defparam \multicast_add_reg[2] .power_up = "low";

dffeas \multicast_add_reg[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[3]~q ),
	.prn(vcc));
defparam \multicast_add_reg[3] .is_wysiwyg = "true";
defparam \multicast_add_reg[3] .power_up = "low";

dffeas \multicast_add_reg[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[4]~q ),
	.prn(vcc));
defparam \multicast_add_reg[4] .is_wysiwyg = "true";
defparam \multicast_add_reg[4] .power_up = "low";

dffeas \multicast_add_reg[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[5]~q ),
	.prn(vcc));
defparam \multicast_add_reg[5] .is_wysiwyg = "true";
defparam \multicast_add_reg[5] .power_up = "low";

dffeas \multicast_add_reg[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[6]~q ),
	.prn(vcc));
defparam \multicast_add_reg[6] .is_wysiwyg = "true";
defparam \multicast_add_reg[6] .power_up = "low";

dffeas \multicast_add_reg[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[7]~q ),
	.prn(vcc));
defparam \multicast_add_reg[7] .is_wysiwyg = "true";
defparam \multicast_add_reg[7] .power_up = "low";

dffeas \multicast_add_reg[8] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[8]~q ),
	.prn(vcc));
defparam \multicast_add_reg[8] .is_wysiwyg = "true";
defparam \multicast_add_reg[8] .power_up = "low";

dffeas \multicast_add_reg[9] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[9]~q ),
	.prn(vcc));
defparam \multicast_add_reg[9] .is_wysiwyg = "true";
defparam \multicast_add_reg[9] .power_up = "low";

dffeas \multicast_add_reg[10] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[10]~q ),
	.prn(vcc));
defparam \multicast_add_reg[10] .is_wysiwyg = "true";
defparam \multicast_add_reg[10] .power_up = "low";

dffeas \multicast_add_reg[11] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[11]~q ),
	.prn(vcc));
defparam \multicast_add_reg[11] .is_wysiwyg = "true";
defparam \multicast_add_reg[11] .power_up = "low";

dffeas \multicast_add_reg[12] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[12]~q ),
	.prn(vcc));
defparam \multicast_add_reg[12] .is_wysiwyg = "true";
defparam \multicast_add_reg[12] .power_up = "low";

dffeas \multicast_add_reg[13] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[13]~q ),
	.prn(vcc));
defparam \multicast_add_reg[13] .is_wysiwyg = "true";
defparam \multicast_add_reg[13] .power_up = "low";

dffeas \multicast_add_reg[14] (
	.clk(mac_rx_clock_connection_clk),
	.d(\multicast_add_reg[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\multicast_add_reg[14]~q ),
	.prn(vcc));
defparam \multicast_add_reg[14] .is_wysiwyg = "true";
defparam \multicast_add_reg[14] .power_up = "low";

cyclonev_lcell_comb \rx_mcast~0 (
	.dataa(!\start_wr_fifo~q ),
	.datab(!\fifo_wr_wait~q ),
	.datac(!\broad_add_reg~q ),
	.datad(!\multicast_add_reg[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_mcast~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_mcast~0 .extended_lut = "off";
defparam \rx_mcast~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \rx_mcast~0 .shared_arith = "off";

cyclonev_lcell_comb \rx_mcast~1 (
	.dataa(!\start_wr_fifo~q ),
	.datab(!\fifo_wr_wait~q ),
	.datac(!\broad_add_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rx_mcast~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rx_mcast~1 .extended_lut = "off";
defparam \rx_mcast~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \rx_mcast~1 .shared_arith = "off";

cyclonev_lcell_comb \always20~6 (
	.dataa(!\start_wr_fifo~q ),
	.datab(!\fifo_wr_wait~q ),
	.datac(!\fifo_wr~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always20~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always20~6 .extended_lut = "off";
defparam \always20~6 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \always20~6 .shared_arith = "off";

cyclonev_lcell_comb \cmd_rcv~0 (
	.dataa(!\sleep_mode_ena~q ),
	.datab(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cmd_rcv~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cmd_rcv~0 .extended_lut = "off";
defparam \cmd_rcv~0 .lut_mask = 64'h7777777777777777;
defparam \cmd_rcv~0 .shared_arith = "off";

cyclonev_lcell_comb \always25~0 (
	.dataa(!\rx_en_s[7]~q ),
	.datab(!\rx_en_s[6]~q ),
	.datac(!\rx_en_s[5]~q ),
	.datad(!\rx_en_s[4]~q ),
	.datae(!\rx_en_s[3]~q ),
	.dataf(!\rx_en_s[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~0 .extended_lut = "off";
defparam \always25~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \always25~0 .shared_arith = "off";

cyclonev_lcell_comb \always25~1 (
	.dataa(!\rx_stat_wren_s[9]~q ),
	.datab(!\rx_stat_wren_s[8]~q ),
	.datac(!\rx_stat_wren_s[11]~q ),
	.datad(!\rx_stat_wren_s[10]~q ),
	.datae(!\rx_en_s[1]~q ),
	.dataf(!\rx_en_s[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~1 .extended_lut = "off";
defparam \always25~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \always25~1 .shared_arith = "off";

cyclonev_lcell_comb \always25~2 (
	.dataa(!\rx_stat_wren_s[2]~q ),
	.datab(!\rx_stat_wren_s[7]~q ),
	.datac(!\rx_stat_wren_s[6]~q ),
	.datad(!\rx_stat_wren_s[5]~q ),
	.datae(!\rx_stat_wren_s[4]~q ),
	.dataf(!\rx_stat_wren_s[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~2 .extended_lut = "off";
defparam \always25~2 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \always25~2 .shared_arith = "off";

cyclonev_lcell_comb \always25~3 (
	.dataa(!\rx_en_s[24]~q ),
	.datab(!\rx_en_s[23]~q ),
	.datac(!\rx_en_s[25]~q ),
	.datad(!\rx_en_s[22]~q ),
	.datae(!\rx_en_s[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~3 .extended_lut = "off";
defparam \always25~3 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always25~3 .shared_arith = "off";

cyclonev_lcell_comb \always25~4 (
	.dataa(!\rx_en_s[19]~q ),
	.datab(!\rx_en_s[18]~q ),
	.datac(!\rx_en_s[17]~q ),
	.datad(!\rx_en_s[16]~q ),
	.datae(!\rx_en_s[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~4 .extended_lut = "off";
defparam \always25~4 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always25~4 .shared_arith = "off";

cyclonev_lcell_comb \always25~5 (
	.dataa(!\rx_en_s[12]~q ),
	.datab(!\rx_en_s[11]~q ),
	.datac(!\rx_en_s[10]~q ),
	.datad(!\rx_en_s[13]~q ),
	.datae(!\rx_en_s[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~5 .extended_lut = "off";
defparam \always25~5 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always25~5 .shared_arith = "off";

cyclonev_lcell_comb \always25~6 (
	.dataa(!\rx_en_s[14]~q ),
	.datab(!\rx_en_s[20]~q ),
	.datac(!\rx_en_s[8]~q ),
	.datad(!\always25~3_combout ),
	.datae(!\always25~4_combout ),
	.dataf(!\always25~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~6 .extended_lut = "off";
defparam \always25~6 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \always25~6 .shared_arith = "off";

cyclonev_lcell_comb \always25~7 (
	.dataa(!\rx_stat_wren_s[1]~q ),
	.datab(!\rx_stat_wren_s[0]~q ),
	.datac(!\always25~0_combout ),
	.datad(!\always25~1_combout ),
	.datae(!\always25~2_combout ),
	.dataf(!\always25~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always25~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always25~7 .extended_lut = "off";
defparam \always25~7 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \always25~7 .shared_arith = "off";

dffeas \rxd_25[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[3]~q ),
	.prn(vcc));
defparam \rxd_25[3] .is_wysiwyg = "true";
defparam \rxd_25[3] .power_up = "low";

dffeas \rxd_25[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[2]~q ),
	.prn(vcc));
defparam \rxd_25[2] .is_wysiwyg = "true";
defparam \rxd_25[2] .power_up = "low";

dffeas \rxd_25[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[1]~q ),
	.prn(vcc));
defparam \rxd_25[1] .is_wysiwyg = "true";
defparam \rxd_25[1] .power_up = "low";

dffeas \rxd_25[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[0]~q ),
	.prn(vcc));
defparam \rxd_25[0] .is_wysiwyg = "true";
defparam \rxd_25[0] .power_up = "low";

dffeas \rxd_25[7] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[7]~q ),
	.prn(vcc));
defparam \rxd_25[7] .is_wysiwyg = "true";
defparam \rxd_25[7] .power_up = "low";

dffeas \rxd_25[6] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[6]~q ),
	.prn(vcc));
defparam \rxd_25[6] .is_wysiwyg = "true";
defparam \rxd_25[6] .power_up = "low";

dffeas \rxd_25[5] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[5]~q ),
	.prn(vcc));
defparam \rxd_25[5] .is_wysiwyg = "true";
defparam \rxd_25[5] .power_up = "low";

dffeas \rxd_25[4] (
	.clk(mac_rx_clock_connection_clk),
	.d(\U_SHIFTTAPS|shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3~portbdataout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\rxd_25[4]~q ),
	.prn(vcc));
defparam \rxd_25[4] .is_wysiwyg = "true";
defparam \rxd_25[4] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_114 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_118 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_115 (
	altera_tse_reset_synchronizer_chain_out,
	ethernet_mode,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
input 	ethernet_mode;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_114 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.din(ethernet_mode),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_114 (
	reset_n,
	din,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_116 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_115 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_115 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_118 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
input 	dreg_1;
output 	dreg_11;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_117 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.din(dreg_1),
	.dreg_1(dreg_11),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_117 (
	reset_n,
	din,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	din;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_118 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_119 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_119 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_119 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_120 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	sleep_ena,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	sleep_ena;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_120 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(sleep_ena),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_120 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_121 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_121 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_121 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_123 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_123 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_123 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_124 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_124 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_124 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_126 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_126 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_126 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_127 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_127 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_rx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_127 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_altshifttaps (
	ram_block5a4,
	ram_block5a5,
	ram_block5a6,
	ram_block5a7,
	ram_block5a0,
	ram_block5a1,
	ram_block5a2,
	ram_block5a3,
	rxclk_ena,
	rxd_8_0,
	rxd_8_1,
	rxd_8_2,
	rxd_8_3,
	rxd_8_4,
	rxd_8_5,
	rxd_8_6,
	rxd_8_7,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	ram_block5a4;
output 	ram_block5a5;
output 	ram_block5a6;
output 	ram_block5a7;
output 	ram_block5a0;
output 	ram_block5a1;
output 	ram_block5a2;
output 	ram_block5a3;
input 	rxclk_ena;
input 	rxd_8_0;
input 	rxd_8_1;
input 	rxd_8_2;
input 	rxd_8_3;
input 	rxd_8_4;
input 	rxd_8_5;
input 	rxd_8_6;
input 	rxd_8_7;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \shift_reg_rtl_0|auto_generated|op_1~1_sumout ;
wire \shift_reg_rtl_0|auto_generated|dffe3a[0]~q ;
wire \shift_reg_rtl_0|auto_generated|op_1~2 ;
wire \shift_reg_rtl_0|auto_generated|op_1~5_sumout ;
wire \shift_reg_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \shift_reg_rtl_0|auto_generated|dffe3a[1]~q ;
wire \shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \shift_reg_rtl_0|auto_generated|op_1~6 ;
wire \shift_reg_rtl_0|auto_generated|op_1~9_sumout ;
wire \shift_reg_rtl_0|auto_generated|dffe3a[2]~q ;
wire \shift_reg_rtl_0|auto_generated|op_1~10 ;
wire \shift_reg_rtl_0|auto_generated|op_1~13_sumout ;
wire \shift_reg_rtl_0|auto_generated|dffe3a[3]~q ;

wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2_PORTBDATAOUT_bus ;
wire [143:0] \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3_PORTBDATAOUT_bus ;

assign ram_block5a4 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4_PORTBDATAOUT_bus [0];

assign ram_block5a5 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5_PORTBDATAOUT_bus [0];

assign ram_block5a6 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6_PORTBDATAOUT_bus [0];

assign ram_block5a7 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7_PORTBDATAOUT_bus [0];

assign ram_block5a0 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0_PORTBDATAOUT_bus [0];

assign ram_block5a1 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1_PORTBDATAOUT_bus [0];

assign ram_block5a2 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2_PORTBDATAOUT_bus [0];

assign ram_block5a3 = \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3_PORTBDATAOUT_bus [0];

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_first_bit_number = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_first_bit_number = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a4 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_first_bit_number = 5;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_first_bit_number = 5;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a5 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_first_bit_number = 6;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_first_bit_number = 6;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a6 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_first_bit_number = 7;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_first_bit_number = 7;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a7 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_first_bit_number = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_first_bit_number = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a0 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_first_bit_number = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_first_bit_number = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a1 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_first_bit_number = 2;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_first_bit_number = 2;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a2 .ram_block_type = "auto";

cyclonev_ram_block \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(mac_rx_clock_connection_clk),
	.clk1(mac_rx_clock_connection_clk),
	.ena0(rxclk_ena),
	.ena1(rxclk_ena),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,rxd_8_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,
\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ,\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\shift_reg_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .clk0_core_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .clk0_input_clock_enable = "ena0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .clk1_output_clock_enable = "ena1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .data_interleave_offset_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .data_interleave_width_in_bits = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_top_1geth:U_GETH|altera_tse_mac_rx:U_RX|altera_tse_altshifttaps:U_SHIFTTAPS|altshift_taps:shift_reg_rtl_0|shift_taps_ffv:auto_generated|altsyncram_1r91:altsyncram4|ALTSYNCRAM";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .mixed_port_feed_through_mode = "dont_care";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .operation_mode = "dual_port";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_data_out_clock = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_first_bit_number = 3;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_address_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_address_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_address_width = 4;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_data_out_clear = "none";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_data_out_clock = "clock1";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_data_width = 1;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_first_address = 0;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_first_bit_number = 3;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_last_address = 15;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_logical_ram_depth = 16;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_logical_ram_width = 8;
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .port_b_read_enable_clock = "clock0";
defparam \shift_reg_rtl_0|auto_generated|altsyncram4|ram_block5a3 .ram_block_type = "auto";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\shift_reg_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|dffe3a[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\shift_reg_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\shift_reg_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\shift_reg_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|dffe3a[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\shift_reg_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \shift_reg_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\shift_reg_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\shift_reg_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|dffe3a[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \shift_reg_rtl_0|auto_generated|op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\shift_reg_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\shift_reg_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\shift_reg_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(),
	.shareout());
defparam \shift_reg_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \shift_reg_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h00000000000000FF;
defparam \shift_reg_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \shift_reg_rtl_0|auto_generated|dffe3a[3] (
	.clk(mac_rx_clock_connection_clk),
	.d(\shift_reg_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\shift_reg_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \shift_reg_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \shift_reg_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_crc328checker (
	altera_tse_reset_synchronizer_chain_out,
	rxclk_ena,
	eof_dly_2,
	frm_type_ok_s_0,
	crc_ok1,
	rxd_25_3,
	rxd_25_2,
	rxd_25_1,
	rxd_25_0,
	rxd_25_7,
	rxd_25_6,
	rxd_25_5,
	rxd_25_4,
	eof,
	mac_rx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
input 	rxclk_ena;
output 	eof_dly_2;
input 	frm_type_ok_s_0;
output 	crc_ok1;
input 	rxd_25_3;
input 	rxd_25_2;
input 	rxd_25_1;
input 	rxd_25_0;
input 	rxd_25_7;
input 	rxd_25_6;
input 	rxd_25_5;
input 	rxd_25_4;
input 	eof;
input 	mac_rx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_GALS|reg_out[7]~q ;
wire \U_GALS|reg_out[9]~q ;
wire \U_GALS|reg_out[11]~q ;
wire \U_GALS|reg_out[24]~q ;
wire \U_GALS|reg_out[3]~q ;
wire \U_GALS|reg_out[2]~q ;
wire \U_GALS|reg_out[16]~q ;
wire \U_GALS|reg_out[0]~q ;
wire \U_GALS|reg_out[4]~q ;
wire \U_GALS|reg_out[19]~q ;
wire \U_GALS|reg_out[20]~q ;
wire \U_GALS|reg_out[29]~q ;
wire \U_GALS|reg_out[22]~q ;
wire \U_GALS|reg_out[27]~q ;
wire \U_GALS|reg_out[23]~q ;
wire \U_GALS|reg_out[26]~q ;
wire \U_GALS|reg_out[30]~q ;
wire \U_GALS|reg_out[31]~q ;
wire \U_GALS|reg_out[28]~q ;
wire \U_GALS|reg_out[25]~q ;
wire \U_GALS|reg_out[21]~q ;
wire \U_GALS|reg_out[18]~q ;
wire \U_GALS|reg_out[17]~q ;
wire \U_GALS|reg_out[15]~q ;
wire \U_GALS|reg_out[14]~q ;
wire \U_GALS|reg_out[13]~q ;
wire \U_GALS|reg_out[12]~q ;
wire \U_GALS|reg_out[10]~q ;
wire \U_GALS|reg_out[8]~q ;
wire \U_GALS|reg_out[6]~q ;
wire \U_GALS|reg_out[5]~q ;
wire \U_GALS|reg_out[1]~q ;
wire \eof_dly[0]~q ;
wire \eof_dly[1]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \Equal0~4_combout ;
wire \Equal0~5_combout ;
wire \Equal0~6_combout ;


IoTOctopus_QSYS_altera_tse_crc32galois8 U_GALS(
	.reg_out_7(\U_GALS|reg_out[7]~q ),
	.reg_out_9(\U_GALS|reg_out[9]~q ),
	.reg_out_11(\U_GALS|reg_out[11]~q ),
	.reg_out_24(\U_GALS|reg_out[24]~q ),
	.reg_out_3(\U_GALS|reg_out[3]~q ),
	.reg_out_2(\U_GALS|reg_out[2]~q ),
	.reg_out_16(\U_GALS|reg_out[16]~q ),
	.reg_out_0(\U_GALS|reg_out[0]~q ),
	.reg_out_4(\U_GALS|reg_out[4]~q ),
	.reg_out_19(\U_GALS|reg_out[19]~q ),
	.reg_out_20(\U_GALS|reg_out[20]~q ),
	.reg_out_29(\U_GALS|reg_out[29]~q ),
	.reg_out_22(\U_GALS|reg_out[22]~q ),
	.reg_out_27(\U_GALS|reg_out[27]~q ),
	.reg_out_23(\U_GALS|reg_out[23]~q ),
	.reg_out_26(\U_GALS|reg_out[26]~q ),
	.reg_out_30(\U_GALS|reg_out[30]~q ),
	.reg_out_31(\U_GALS|reg_out[31]~q ),
	.reg_out_28(\U_GALS|reg_out[28]~q ),
	.reg_out_25(\U_GALS|reg_out[25]~q ),
	.reg_out_21(\U_GALS|reg_out[21]~q ),
	.reg_out_18(\U_GALS|reg_out[18]~q ),
	.reg_out_17(\U_GALS|reg_out[17]~q ),
	.reg_out_15(\U_GALS|reg_out[15]~q ),
	.reg_out_14(\U_GALS|reg_out[14]~q ),
	.reg_out_13(\U_GALS|reg_out[13]~q ),
	.reg_out_12(\U_GALS|reg_out[12]~q ),
	.reg_out_10(\U_GALS|reg_out[10]~q ),
	.reg_out_8(\U_GALS|reg_out[8]~q ),
	.reg_out_6(\U_GALS|reg_out[6]~q ),
	.reg_out_5(\U_GALS|reg_out[5]~q ),
	.reg_out_1(\U_GALS|reg_out[1]~q ),
	.rst(altera_tse_reset_synchronizer_chain_out),
	.clk_ena(rxclk_ena),
	.frm_type_ok_s_0(frm_type_ok_s_0),
	.rxd_25_3(rxd_25_3),
	.rxd_25_2(rxd_25_2),
	.rxd_25_1(rxd_25_1),
	.rxd_25_0(rxd_25_0),
	.rxd_25_7(rxd_25_7),
	.rxd_25_6(rxd_25_6),
	.rxd_25_5(rxd_25_5),
	.rxd_25_4(rxd_25_4),
	.clk(mac_rx_clock_connection_clk));

dffeas \eof_dly[2] (
	.clk(mac_rx_clock_connection_clk),
	.d(\eof_dly[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(eof_dly_2),
	.prn(vcc));
defparam \eof_dly[2] .is_wysiwyg = "true";
defparam \eof_dly[2] .power_up = "low";

dffeas crc_ok(
	.clk(mac_rx_clock_connection_clk),
	.d(\Equal0~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(crc_ok1),
	.prn(vcc));
defparam crc_ok.is_wysiwyg = "true";
defparam crc_ok.power_up = "low";

dffeas \eof_dly[0] (
	.clk(mac_rx_clock_connection_clk),
	.d(eof),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\eof_dly[0]~q ),
	.prn(vcc));
defparam \eof_dly[0] .is_wysiwyg = "true";
defparam \eof_dly[0] .power_up = "low";

dffeas \eof_dly[1] (
	.clk(mac_rx_clock_connection_clk),
	.d(\eof_dly[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(rxclk_ena),
	.q(\eof_dly[1]~q ),
	.prn(vcc));
defparam \eof_dly[1] .is_wysiwyg = "true";
defparam \eof_dly[1] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\U_GALS|reg_out[7]~q ),
	.datab(!\U_GALS|reg_out[9]~q ),
	.datac(!\U_GALS|reg_out[11]~q ),
	.datad(!\U_GALS|reg_out[24]~q ),
	.datae(!\U_GALS|reg_out[3]~q ),
	.dataf(!\U_GALS|reg_out[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\U_GALS|reg_out[16]~q ),
	.datab(!\U_GALS|reg_out[0]~q ),
	.datac(!\U_GALS|reg_out[4]~q ),
	.datad(!\U_GALS|reg_out[19]~q ),
	.datae(!\U_GALS|reg_out[20]~q ),
	.dataf(!\U_GALS|reg_out[29]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\U_GALS|reg_out[22]~q ),
	.datab(!\U_GALS|reg_out[27]~q ),
	.datac(!\U_GALS|reg_out[23]~q ),
	.datad(!\U_GALS|reg_out[26]~q ),
	.datae(!\U_GALS|reg_out[30]~q ),
	.dataf(!\U_GALS|reg_out[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!\U_GALS|reg_out[28]~q ),
	.datab(!\U_GALS|reg_out[25]~q ),
	.datac(!\U_GALS|reg_out[21]~q ),
	.datad(!\U_GALS|reg_out[18]~q ),
	.datae(!\U_GALS|reg_out[17]~q ),
	.dataf(!\U_GALS|reg_out[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!\U_GALS|reg_out[14]~q ),
	.datab(!\U_GALS|reg_out[13]~q ),
	.datac(!\U_GALS|reg_out[12]~q ),
	.datad(!\U_GALS|reg_out[10]~q ),
	.datae(!\U_GALS|reg_out[8]~q ),
	.dataf(!\U_GALS|reg_out[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~5 (
	.dataa(!\U_GALS|reg_out[5]~q ),
	.datab(!\U_GALS|reg_out[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'h7777777777777777;
defparam \Equal0~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~6 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~1_combout ),
	.datac(!\Equal0~2_combout ),
	.datad(!\Equal0~3_combout ),
	.datae(!\Equal0~4_combout ),
	.dataf(!\Equal0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~6 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_crc32galois8 (
	reg_out_7,
	reg_out_9,
	reg_out_11,
	reg_out_24,
	reg_out_3,
	reg_out_2,
	reg_out_16,
	reg_out_0,
	reg_out_4,
	reg_out_19,
	reg_out_20,
	reg_out_29,
	reg_out_22,
	reg_out_27,
	reg_out_23,
	reg_out_26,
	reg_out_30,
	reg_out_31,
	reg_out_28,
	reg_out_25,
	reg_out_21,
	reg_out_18,
	reg_out_17,
	reg_out_15,
	reg_out_14,
	reg_out_13,
	reg_out_12,
	reg_out_10,
	reg_out_8,
	reg_out_6,
	reg_out_5,
	reg_out_1,
	rst,
	clk_ena,
	frm_type_ok_s_0,
	rxd_25_3,
	rxd_25_2,
	rxd_25_1,
	rxd_25_0,
	rxd_25_7,
	rxd_25_6,
	rxd_25_5,
	rxd_25_4,
	clk)/* synthesis synthesis_greybox=1 */;
output 	reg_out_7;
output 	reg_out_9;
output 	reg_out_11;
output 	reg_out_24;
output 	reg_out_3;
output 	reg_out_2;
output 	reg_out_16;
output 	reg_out_0;
output 	reg_out_4;
output 	reg_out_19;
output 	reg_out_20;
output 	reg_out_29;
output 	reg_out_22;
output 	reg_out_27;
output 	reg_out_23;
output 	reg_out_26;
output 	reg_out_30;
output 	reg_out_31;
output 	reg_out_28;
output 	reg_out_25;
output 	reg_out_21;
output 	reg_out_18;
output 	reg_out_17;
output 	reg_out_15;
output 	reg_out_14;
output 	reg_out_13;
output 	reg_out_12;
output 	reg_out_10;
output 	reg_out_8;
output 	reg_out_6;
output 	reg_out_5;
output 	reg_out_1;
input 	rst;
input 	clk_ena;
input 	frm_type_ok_s_0;
input 	rxd_25_3;
input 	rxd_25_2;
input 	rxd_25_1;
input 	rxd_25_0;
input 	rxd_25_7;
input 	rxd_25_6;
input 	rxd_25_5;
input 	rxd_25_4;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \o[7]~combout ;
wire \o[9]~combout ;
wire \o[11]~combout ;
wire \o[24]~combout ;
wire \o[3]~combout ;
wire \o[2]~combout ;
wire \o[16]~combout ;
wire \o[0]~combout ;
wire \o[4]~combout ;
wire \o[19]~0_combout ;
wire \o[19]~combout ;
wire \o[20]~combout ;
wire \o[29]~combout ;
wire \o[22]~combout ;
wire \o[27]~combout ;
wire \o[23]~combout ;
wire \o1[0]~combout ;
wire \o[26]~combout ;
wire \o[30]~combout ;
wire \o[31]~combout ;
wire \o[28]~combout ;
wire \o[25]~combout ;
wire \o[21]~combout ;
wire \o[18]~1_combout ;
wire \o[18]~combout ;
wire \o[17]~combout ;
wire \o[15]~combout ;
wire \o[14]~combout ;
wire \o[13]~combout ;
wire \o[12]~combout ;
wire \o[10]~combout ;
wire \o[8]~combout ;
wire \o[6]~combout ;
wire \o[5]~combout ;
wire \o[1]~combout ;


dffeas \reg_out[7] (
	.clk(clk),
	.d(\o[7]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_7),
	.prn(vcc));
defparam \reg_out[7] .is_wysiwyg = "true";
defparam \reg_out[7] .power_up = "low";

dffeas \reg_out[9] (
	.clk(clk),
	.d(\o[9]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_9),
	.prn(vcc));
defparam \reg_out[9] .is_wysiwyg = "true";
defparam \reg_out[9] .power_up = "low";

dffeas \reg_out[11] (
	.clk(clk),
	.d(\o[11]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_11),
	.prn(vcc));
defparam \reg_out[11] .is_wysiwyg = "true";
defparam \reg_out[11] .power_up = "low";

dffeas \reg_out[24] (
	.clk(clk),
	.d(\o[24]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_24),
	.prn(vcc));
defparam \reg_out[24] .is_wysiwyg = "true";
defparam \reg_out[24] .power_up = "low";

dffeas \reg_out[3] (
	.clk(clk),
	.d(\o[3]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_3),
	.prn(vcc));
defparam \reg_out[3] .is_wysiwyg = "true";
defparam \reg_out[3] .power_up = "low";

dffeas \reg_out[2] (
	.clk(clk),
	.d(\o[2]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_2),
	.prn(vcc));
defparam \reg_out[2] .is_wysiwyg = "true";
defparam \reg_out[2] .power_up = "low";

dffeas \reg_out[16] (
	.clk(clk),
	.d(\o[16]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_16),
	.prn(vcc));
defparam \reg_out[16] .is_wysiwyg = "true";
defparam \reg_out[16] .power_up = "low";

dffeas \reg_out[0] (
	.clk(clk),
	.d(\o[0]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_0),
	.prn(vcc));
defparam \reg_out[0] .is_wysiwyg = "true";
defparam \reg_out[0] .power_up = "low";

dffeas \reg_out[4] (
	.clk(clk),
	.d(\o[4]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_4),
	.prn(vcc));
defparam \reg_out[4] .is_wysiwyg = "true";
defparam \reg_out[4] .power_up = "low";

dffeas \reg_out[19] (
	.clk(clk),
	.d(\o[19]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_19),
	.prn(vcc));
defparam \reg_out[19] .is_wysiwyg = "true";
defparam \reg_out[19] .power_up = "low";

dffeas \reg_out[20] (
	.clk(clk),
	.d(\o[20]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_20),
	.prn(vcc));
defparam \reg_out[20] .is_wysiwyg = "true";
defparam \reg_out[20] .power_up = "low";

dffeas \reg_out[29] (
	.clk(clk),
	.d(\o[29]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_29),
	.prn(vcc));
defparam \reg_out[29] .is_wysiwyg = "true";
defparam \reg_out[29] .power_up = "low";

dffeas \reg_out[22] (
	.clk(clk),
	.d(\o[22]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_22),
	.prn(vcc));
defparam \reg_out[22] .is_wysiwyg = "true";
defparam \reg_out[22] .power_up = "low";

dffeas \reg_out[27] (
	.clk(clk),
	.d(\o[27]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_27),
	.prn(vcc));
defparam \reg_out[27] .is_wysiwyg = "true";
defparam \reg_out[27] .power_up = "low";

dffeas \reg_out[23] (
	.clk(clk),
	.d(\o[23]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_23),
	.prn(vcc));
defparam \reg_out[23] .is_wysiwyg = "true";
defparam \reg_out[23] .power_up = "low";

dffeas \reg_out[26] (
	.clk(clk),
	.d(\o[26]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_26),
	.prn(vcc));
defparam \reg_out[26] .is_wysiwyg = "true";
defparam \reg_out[26] .power_up = "low";

dffeas \reg_out[30] (
	.clk(clk),
	.d(\o[30]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(frm_type_ok_s_0),
	.sload(gnd),
	.ena(clk_ena),
	.q(reg_out_30),
	.prn(vcc));
defparam \reg_out[30] .is_wysiwyg = "true";
defparam \reg_out[30] .power_up = "low";

dffeas \reg_out[31] (
	.clk(clk),
	.d(\o[31]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_31),
	.prn(vcc));
defparam \reg_out[31] .is_wysiwyg = "true";
defparam \reg_out[31] .power_up = "low";

dffeas \reg_out[28] (
	.clk(clk),
	.d(\o[28]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_28),
	.prn(vcc));
defparam \reg_out[28] .is_wysiwyg = "true";
defparam \reg_out[28] .power_up = "low";

dffeas \reg_out[25] (
	.clk(clk),
	.d(\o[25]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_25),
	.prn(vcc));
defparam \reg_out[25] .is_wysiwyg = "true";
defparam \reg_out[25] .power_up = "low";

dffeas \reg_out[21] (
	.clk(clk),
	.d(\o[21]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_21),
	.prn(vcc));
defparam \reg_out[21] .is_wysiwyg = "true";
defparam \reg_out[21] .power_up = "low";

dffeas \reg_out[18] (
	.clk(clk),
	.d(\o[18]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_18),
	.prn(vcc));
defparam \reg_out[18] .is_wysiwyg = "true";
defparam \reg_out[18] .power_up = "low";

dffeas \reg_out[17] (
	.clk(clk),
	.d(\o[17]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_17),
	.prn(vcc));
defparam \reg_out[17] .is_wysiwyg = "true";
defparam \reg_out[17] .power_up = "low";

dffeas \reg_out[15] (
	.clk(clk),
	.d(\o[15]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_15),
	.prn(vcc));
defparam \reg_out[15] .is_wysiwyg = "true";
defparam \reg_out[15] .power_up = "low";

dffeas \reg_out[14] (
	.clk(clk),
	.d(\o[14]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_14),
	.prn(vcc));
defparam \reg_out[14] .is_wysiwyg = "true";
defparam \reg_out[14] .power_up = "low";

dffeas \reg_out[13] (
	.clk(clk),
	.d(\o[13]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_13),
	.prn(vcc));
defparam \reg_out[13] .is_wysiwyg = "true";
defparam \reg_out[13] .power_up = "low";

dffeas \reg_out[12] (
	.clk(clk),
	.d(\o[12]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_12),
	.prn(vcc));
defparam \reg_out[12] .is_wysiwyg = "true";
defparam \reg_out[12] .power_up = "low";

dffeas \reg_out[10] (
	.clk(clk),
	.d(\o[10]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_10),
	.prn(vcc));
defparam \reg_out[10] .is_wysiwyg = "true";
defparam \reg_out[10] .power_up = "low";

dffeas \reg_out[8] (
	.clk(clk),
	.d(\o[8]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_8),
	.prn(vcc));
defparam \reg_out[8] .is_wysiwyg = "true";
defparam \reg_out[8] .power_up = "low";

dffeas \reg_out[6] (
	.clk(clk),
	.d(\o[6]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_6),
	.prn(vcc));
defparam \reg_out[6] .is_wysiwyg = "true";
defparam \reg_out[6] .power_up = "low";

dffeas \reg_out[5] (
	.clk(clk),
	.d(\o[5]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_5),
	.prn(vcc));
defparam \reg_out[5] .is_wysiwyg = "true";
defparam \reg_out[5] .power_up = "low";

dffeas \reg_out[1] (
	.clk(clk),
	.d(\o[1]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(frm_type_ok_s_0),
	.ena(clk_ena),
	.q(reg_out_1),
	.prn(vcc));
defparam \reg_out[1] .is_wysiwyg = "true";
defparam \reg_out[1] .power_up = "low";

cyclonev_lcell_comb \o[7] (
	.dataa(!reg_out_0),
	.datab(!reg_out_15),
	.datac(!reg_out_6),
	.datad(!reg_out_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[7] .extended_lut = "off";
defparam \o[7] .lut_mask = 64'h6996699669966996;
defparam \o[7] .shared_arith = "off";

cyclonev_lcell_comb \o[9] (
	.dataa(!reg_out_7),
	.datab(!reg_out_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[9] .extended_lut = "off";
defparam \o[9] .lut_mask = 64'h6666666666666666;
defparam \o[9] .shared_arith = "off";

cyclonev_lcell_comb \o[11] (
	.dataa(!reg_out_3),
	.datab(!reg_out_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[11] .extended_lut = "off";
defparam \o[11] .lut_mask = 64'h6666666666666666;
defparam \o[11] .shared_arith = "off";

cyclonev_lcell_comb \o[24] (
	.dataa(!rxd_25_0),
	.datab(!reg_out_7),
	.datac(!reg_out_2),
	.datad(!reg_out_0),
	.datae(!reg_out_4),
	.dataf(!reg_out_5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[24] .extended_lut = "off";
defparam \o[24] .lut_mask = 64'h6996966996696996;
defparam \o[24] .shared_arith = "off";

cyclonev_lcell_comb \o[3] (
	.dataa(!reg_out_11),
	.datab(!reg_out_2),
	.datac(!reg_out_5),
	.datad(!reg_out_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[3] .extended_lut = "off";
defparam \o[3] .lut_mask = 64'h6996699669966996;
defparam \o[3] .shared_arith = "off";

cyclonev_lcell_comb \o[2] (
	.dataa(!reg_out_0),
	.datab(!reg_out_4),
	.datac(!reg_out_10),
	.datad(!reg_out_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[2] .extended_lut = "off";
defparam \o[2] .lut_mask = 64'h6996699669966996;
defparam \o[2] .shared_arith = "off";

cyclonev_lcell_comb \o[16] (
	.dataa(!reg_out_24),
	.datab(!reg_out_3),
	.datac(!reg_out_2),
	.datad(!reg_out_0),
	.datae(!reg_out_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[16] .extended_lut = "off";
defparam \o[16] .lut_mask = 64'h9669699696696996;
defparam \o[16] .shared_arith = "off";

cyclonev_lcell_comb \o[0] (
	.dataa(!reg_out_2),
	.datab(!reg_out_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[0] .extended_lut = "off";
defparam \o[0] .lut_mask = 64'h6666666666666666;
defparam \o[0] .shared_arith = "off";

cyclonev_lcell_comb \o[4] (
	.dataa(!reg_out_3),
	.datab(!reg_out_2),
	.datac(!reg_out_0),
	.datad(!reg_out_12),
	.datae(!reg_out_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[4] .extended_lut = "off";
defparam \o[4] .lut_mask = 64'h9669699696696996;
defparam \o[4] .shared_arith = "off";

cyclonev_lcell_comb \o[19]~0 (
	.dataa(!reg_out_7),
	.datab(!reg_out_3),
	.datac(!reg_out_2),
	.datad(!reg_out_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[19]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[19]~0 .extended_lut = "off";
defparam \o[19]~0 .lut_mask = 64'h6996699669966996;
defparam \o[19]~0 .shared_arith = "off";

cyclonev_lcell_comb \o[19] (
	.dataa(!reg_out_27),
	.datab(!reg_out_6),
	.datac(!reg_out_5),
	.datad(!\o[19]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[19] .extended_lut = "off";
defparam \o[19] .lut_mask = 64'h6996699669966996;
defparam \o[19] .shared_arith = "off";

cyclonev_lcell_comb \o[20] (
	.dataa(!reg_out_7),
	.datab(!reg_out_3),
	.datac(!reg_out_4),
	.datad(!reg_out_28),
	.datae(!reg_out_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[20] .extended_lut = "off";
defparam \o[20] .lut_mask = 64'h9669699696696996;
defparam \o[20] .shared_arith = "off";

cyclonev_lcell_comb \o[29] (
	.dataa(!rxd_25_5),
	.datab(!reg_out_7),
	.datac(!reg_out_0),
	.datad(!reg_out_6),
	.datae(!reg_out_5),
	.dataf(!reg_out_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[29] .extended_lut = "off";
defparam \o[29] .lut_mask = 64'h6996966996696996;
defparam \o[29] .shared_arith = "off";

cyclonev_lcell_comb \o[22] (
	.dataa(!reg_out_3),
	.datab(!reg_out_2),
	.datac(!reg_out_30),
	.datad(!reg_out_6),
	.datae(!reg_out_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[22] .extended_lut = "off";
defparam \o[22] .lut_mask = 64'h9669699696696996;
defparam \o[22] .shared_arith = "off";

cyclonev_lcell_comb \o[27] (
	.dataa(!rxd_25_3),
	.datab(!reg_out_7),
	.datac(!reg_out_3),
	.datad(!reg_out_4),
	.datae(!reg_out_5),
	.dataf(!reg_out_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[27] .extended_lut = "off";
defparam \o[27] .lut_mask = 64'h6996966996696996;
defparam \o[27] .shared_arith = "off";

cyclonev_lcell_comb \o[23] (
	.dataa(!reg_out_7),
	.datab(!reg_out_3),
	.datac(!reg_out_4),
	.datad(!reg_out_31),
	.datae(!reg_out_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[23] .extended_lut = "off";
defparam \o[23] .lut_mask = 64'h9669699696696996;
defparam \o[23] .shared_arith = "off";

cyclonev_lcell_comb \o1[0] (
	.dataa(!reg_out_3),
	.datab(!reg_out_2),
	.datac(!reg_out_0),
	.datad(!reg_out_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o1[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o1[0] .extended_lut = "off";
defparam \o1[0] .lut_mask = 64'h6996699669966996;
defparam \o1[0] .shared_arith = "off";

cyclonev_lcell_comb \o[26] (
	.dataa(!rxd_25_2),
	.datab(!reg_out_7),
	.datac(!reg_out_4),
	.datad(!reg_out_1),
	.datae(!\o1[0]~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[26] .extended_lut = "off";
defparam \o[26] .lut_mask = 64'h9669699696696996;
defparam \o[26] .shared_arith = "off";

cyclonev_lcell_comb \o[30] (
	.dataa(!rxd_25_6),
	.datab(!reg_out_7),
	.datac(!reg_out_0),
	.datad(!reg_out_6),
	.datae(!reg_out_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[30] .extended_lut = "off";
defparam \o[30] .lut_mask = 64'h9669699696696996;
defparam \o[30] .shared_arith = "off";

cyclonev_lcell_comb \o[31] (
	.dataa(!rxd_25_7),
	.datab(!reg_out_7),
	.datac(!reg_out_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[31] .extended_lut = "off";
defparam \o[31] .lut_mask = 64'h9696969696969696;
defparam \o[31] .shared_arith = "off";

cyclonev_lcell_comb \o[28] (
	.dataa(!rxd_25_4),
	.datab(!reg_out_0),
	.datac(!reg_out_4),
	.datad(!reg_out_6),
	.datae(!reg_out_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[28] .extended_lut = "off";
defparam \o[28] .lut_mask = 64'h9669699696696996;
defparam \o[28] .shared_arith = "off";

cyclonev_lcell_comb \o[25] (
	.dataa(!rxd_25_1),
	.datab(!reg_out_5),
	.datac(!reg_out_1),
	.datad(!\o1[0]~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[25] .extended_lut = "off";
defparam \o[25] .lut_mask = 64'h6996699669966996;
defparam \o[25] .shared_arith = "off";

cyclonev_lcell_comb \o[21] (
	.dataa(!reg_out_7),
	.datab(!reg_out_2),
	.datac(!reg_out_4),
	.datad(!reg_out_29),
	.datae(!reg_out_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[21] .extended_lut = "off";
defparam \o[21] .lut_mask = 64'h9669699696696996;
defparam \o[21] .shared_arith = "off";

cyclonev_lcell_comb \o[18]~1 (
	.dataa(!reg_out_2),
	.datab(!reg_out_26),
	.datac(!reg_out_6),
	.datad(!reg_out_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[18]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[18]~1 .extended_lut = "off";
defparam \o[18]~1 .lut_mask = 64'h6996699669966996;
defparam \o[18]~1 .shared_arith = "off";

cyclonev_lcell_comb \o[18] (
	.dataa(!reg_out_0),
	.datab(!reg_out_4),
	.datac(!reg_out_1),
	.datad(!\o[18]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[18] .extended_lut = "off";
defparam \o[18] .lut_mask = 64'h6996699669966996;
defparam \o[18] .shared_arith = "off";

cyclonev_lcell_comb \o[17] (
	.dataa(!reg_out_3),
	.datab(!reg_out_0),
	.datac(!reg_out_4),
	.datad(!reg_out_25),
	.datae(!reg_out_5),
	.dataf(!reg_out_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[17] .extended_lut = "off";
defparam \o[17] .lut_mask = 64'h6996966996696996;
defparam \o[17] .shared_arith = "off";

cyclonev_lcell_comb \o[15] (
	.dataa(!reg_out_7),
	.datab(!reg_out_3),
	.datac(!reg_out_2),
	.datad(!reg_out_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[15] .extended_lut = "off";
defparam \o[15] .lut_mask = 64'h6996699669966996;
defparam \o[15] .shared_arith = "off";

cyclonev_lcell_comb \o[14] (
	.dataa(!reg_out_2),
	.datab(!reg_out_22),
	.datac(!reg_out_6),
	.datad(!reg_out_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[14] .extended_lut = "off";
defparam \o[14] .lut_mask = 64'h6996699669966996;
defparam \o[14] .shared_arith = "off";

cyclonev_lcell_comb \o[13] (
	.dataa(!reg_out_0),
	.datab(!reg_out_21),
	.datac(!reg_out_5),
	.datad(!reg_out_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[13] .extended_lut = "off";
defparam \o[13] .lut_mask = 64'h6996699669966996;
defparam \o[13] .shared_arith = "off";

cyclonev_lcell_comb \o[12] (
	.dataa(!reg_out_0),
	.datab(!reg_out_4),
	.datac(!reg_out_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[12] .extended_lut = "off";
defparam \o[12] .lut_mask = 64'h9696969696969696;
defparam \o[12] .shared_arith = "off";

cyclonev_lcell_comb \o[10] (
	.dataa(!reg_out_2),
	.datab(!reg_out_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[10] .extended_lut = "off";
defparam \o[10] .lut_mask = 64'h6666666666666666;
defparam \o[10] .shared_arith = "off";

cyclonev_lcell_comb \o[8] (
	.dataa(!reg_out_7),
	.datab(!reg_out_16),
	.datac(!reg_out_6),
	.datad(!reg_out_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[8] .extended_lut = "off";
defparam \o[8] .lut_mask = 64'h6996699669966996;
defparam \o[8] .shared_arith = "off";

cyclonev_lcell_comb \o[6] (
	.dataa(!reg_out_4),
	.datab(!reg_out_14),
	.datac(!reg_out_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[6] .extended_lut = "off";
defparam \o[6] .lut_mask = 64'h9696969696969696;
defparam \o[6] .shared_arith = "off";

cyclonev_lcell_comb \o[5] (
	.dataa(!reg_out_7),
	.datab(!reg_out_3),
	.datac(!reg_out_4),
	.datad(!reg_out_13),
	.datae(!reg_out_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[5] .extended_lut = "off";
defparam \o[5] .lut_mask = 64'h9669699696696996;
defparam \o[5] .shared_arith = "off";

cyclonev_lcell_comb \o[1] (
	.dataa(!reg_out_9),
	.datab(!reg_out_3),
	.datac(!reg_out_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[1] .extended_lut = "off";
defparam \o[1] .lut_mask = 64'h9696969696969696;
defparam \o[1] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_mac_tx (
	q_b_9,
	eop_sft_0,
	q_b_8,
	q_b_4,
	dout_reg_sft_28,
	q_b_0,
	dout_reg_sft_24,
	q_b_5,
	dout_reg_sft_29,
	q_b_1,
	dout_reg_sft_25,
	q_b_6,
	dout_reg_sft_30,
	q_b_2,
	dout_reg_sft_26,
	q_b_7,
	dout_reg_sft_31,
	q_b_3,
	dout_reg_sft_27,
	tx_ff_uflow1,
	txclk_ena,
	altera_tse_reset_synchronizer_chain_out,
	tx_empty,
	tx_data_int_7,
	dreg_1,
	tx_en_s_1,
	rd_14_4,
	rd_14_0,
	rd_14_5,
	rd_14_1,
	rd_14_6,
	rd_14_2,
	rd_14_7,
	rd_14_3,
	tx_err1,
	tx_eop_int,
	empty_flag,
	always9,
	col_int1,
	always91,
	tx_rden_mii1,
	tx_rden_int,
	always92,
	mac_ena,
	tx_sav_int,
	ethernet_mode,
	dreg_11,
	tx_stat_1,
	sop_reg,
	tx_stat_rden1,
	sleep_ena,
	dreg_12,
	m_rx_crs,
	tx_stat_0,
	GND_port,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	q_b_9;
input 	eop_sft_0;
input 	q_b_8;
input 	q_b_4;
input 	dout_reg_sft_28;
input 	q_b_0;
input 	dout_reg_sft_24;
input 	q_b_5;
input 	dout_reg_sft_29;
input 	q_b_1;
input 	dout_reg_sft_25;
input 	q_b_6;
input 	dout_reg_sft_30;
input 	q_b_2;
input 	dout_reg_sft_26;
input 	q_b_7;
input 	dout_reg_sft_31;
input 	q_b_3;
input 	dout_reg_sft_27;
output 	tx_ff_uflow1;
input 	txclk_ena;
input 	altera_tse_reset_synchronizer_chain_out;
input 	tx_empty;
input 	tx_data_int_7;
output 	dreg_1;
output 	tx_en_s_1;
output 	rd_14_4;
output 	rd_14_0;
output 	rd_14_5;
output 	rd_14_1;
output 	rd_14_6;
output 	rd_14_2;
output 	rd_14_7;
output 	rd_14_3;
output 	tx_err1;
input 	tx_eop_int;
input 	empty_flag;
output 	always9;
output 	col_int1;
output 	always91;
output 	tx_rden_mii1;
output 	tx_rden_int;
output 	always92;
input 	mac_ena;
input 	tx_sav_int;
input 	ethernet_mode;
output 	dreg_11;
input 	tx_stat_1;
input 	sop_reg;
output 	tx_stat_rden1;
input 	sleep_ena;
input 	dreg_12;
input 	m_rx_crs;
input 	tx_stat_0;
input 	GND_port;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_4|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_7|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_MAGIC_ENA|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_SLEEP_ENA|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \gm_rx_col_reg~q ;
wire \gm_rx_col_reg~0_combout ;
wire \U_CRC|U_CTL|eof_dly[5]~q ;
wire \U_CRC|U_GALS|reg_out[0]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[10]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[11]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[12]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[13]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[14]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[15]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[16]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[17]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[18]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[19]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[1]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[20]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[21]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[22]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[23]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[24]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[25]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[26]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[27]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[28]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[29]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[2]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[30]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[31]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[3]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[4]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[5]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[6]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[7]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[8]~_wirecell_combout ;
wire \U_CRC|U_GALS|reg_out[9]~_wirecell_combout ;
wire \gm_rx_col_reg2~q ;
wire \always3~0_combout ;
wire \always9~0_combout ;
wire \eop_0~1_combout ;
wire \always9~2_combout ;
wire \tx_rden~q ;
wire \tx_rden_d1~q ;
wire \eop_0~0_combout ;
wire \frm_rd~0_combout ;
wire \frm_rd[0]~q ;
wire \eop_0~2_combout ;
wire \always6~0_combout ;
wire \frm_rd[2]~q ;
wire \tx_ff_uflow~0_combout ;
wire \frm_cnt[0]~3_combout ;
wire \frm_cnt[2]~7_combout ;
wire \frm_cnt[2]~q ;
wire \frm_cnt[3]~6_combout ;
wire \frm_cnt[3]~q ;
wire \Add0~0_combout ;
wire \frm_cnt[4]~5_combout ;
wire \frm_cnt[4]~q ;
wire \frm_cnt[5]~4_combout ;
wire \frm_cnt[5]~q ;
wire \Equal0~0_combout ;
wire \frm_cnt[1]~0_combout ;
wire \frm_cnt[4]~1_combout ;
wire \frm_cnt[0]~8_combout ;
wire \frm_cnt[0]~q ;
wire \always6~2_combout ;
wire \frm_cnt[1]~2_combout ;
wire \frm_cnt[1]~q ;
wire \LessThan0~0_combout ;
wire \always6~1_combout ;
wire \frm_rd[1]~q ;
wire \always7~0_combout ;
wire \pad_cnt[5]~0_combout ;
wire \Add1~0_combout ;
wire \pad_cnt[2]~5_combout ;
wire \pad_cnt[2]~q ;
wire \Add1~1_combout ;
wire \pad_cnt[3]~4_combout ;
wire \pad_cnt[3]~q ;
wire \pad_cnt[4]~6_combout ;
wire \pad_cnt[4]~q ;
wire \Add1~2_combout ;
wire \pad_cnt[5]~3_combout ;
wire \pad_cnt[5]~q ;
wire \Equal3~0_combout ;
wire \Equal1~0_combout ;
wire \always7~1_combout ;
wire \pad_cnt~2_combout ;
wire \pad_cnt[0]~q ;
wire \pad_cnt[1]~1_combout ;
wire \pad_cnt[1]~q ;
wire \pad_wait~0_combout ;
wire \pad_wait~q ;
wire \tx_ipg_len_int~0_combout ;
wire \tx_ipg_len_int[0]~q ;
wire \tx_ipg_len_int~1_combout ;
wire \tx_ipg_len_int[1]~q ;
wire \gap_cnt~1_combout ;
wire \gap_cnt[1]~q ;
wire \tx_ipg_len_int~3_combout ;
wire \tx_ipg_len_int[3]~q ;
wire \tx_ipg_len_int~2_combout ;
wire \tx_ipg_len_int[2]~q ;
wire \Add2~1_combout ;
wire \gap_cnt~3_combout ;
wire \gap_cnt[2]~q ;
wire \Add2~2_combout ;
wire \gap_cnt~4_combout ;
wire \gap_cnt[3]~q ;
wire \tx_ipg_len_int~4_combout ;
wire \tx_ipg_len_int[4]~q ;
wire \Add2~0_combout ;
wire \gap_cnt~2_combout ;
wire \gap_cnt[4]~q ;
wire \Equal6~0_combout ;
wire \always13~9_combout ;
wire \always13~10_combout ;
wire \Add4~0_combout ;
wire \always13~11_combout ;
wire \always13~3_combout ;
wire \gap_12_b~q ;
wire \always13~8_combout ;
wire \gap_run[3]~q ;
wire \always13~2_combout ;
wire \gap_run[4]~q ;
wire \gap_cnt~0_combout ;
wire \gap_cnt[0]~q ;
wire \always13~5_combout ;
wire \always13~6_combout ;
wire \gap_12~q ;
wire \always13~7_combout ;
wire \gap_run[0]~q ;
wire \always13~4_combout ;
wire \gap_run[1]~q ;
wire \always13~1_combout ;
wire \gap_run[2]~q ;
wire \always13~0_combout ;
wire \gap_wait~q ;
wire \crc_fwd~0_combout ;
wire \crc_fwd~q ;
wire \always17~0_combout ;
wire \eop~13_combout ;
wire \eop[1]~q ;
wire \eop~15_combout ;
wire \eop[2]~q ;
wire \eop~14_combout ;
wire \eop[3]~q ;
wire \eop[4]~q ;
wire \eop~12_combout ;
wire \eop[5]~q ;
wire \eop~11_combout ;
wire \eop[6]~q ;
wire \eop~10_combout ;
wire \eop[7]~q ;
wire \eop~9_combout ;
wire \eop[8]~q ;
wire \eop~8_combout ;
wire \eop[9]~q ;
wire \eop~6_combout ;
wire \eop[10]~q ;
wire \eop~4_combout ;
wire \eop[11]~q ;
wire \eop~2_combout ;
wire \eop[12]~q ;
wire \eop~0_combout ;
wire \eop[13]~q ;
wire \eop~7_combout ;
wire \eop[14]~q ;
wire \eop~5_combout ;
wire \eop[15]~q ;
wire \eop~3_combout ;
wire \eop[16]~q ;
wire \eop~1_combout ;
wire \eop[17]~q ;
wire \tx_en_s~2_combout ;
wire \sop~0_combout ;
wire \sop[1]~q ;
wire \sop[2]~q ;
wire \sop[3]~q ;
wire \sop[4]~q ;
wire \tx_en_s[0]~q ;
wire \preamb_cnt~2_combout ;
wire \preamb_cnt[0]~q ;
wire \preamb_cnt~1_combout ;
wire \preamb_cnt[1]~q ;
wire \preamb_cnt~0_combout ;
wire \preamb_cnt[2]~q ;
wire \always19~3_combout ;
wire \preamb_run[0]~q ;
wire \always19~4_combout ;
wire \preamb_run[1]~q ;
wire \always19~2_combout ;
wire \preamb_run[2]~q ;
wire \always19~1_combout ;
wire \preamb_wait~0_combout ;
wire \preamb_wait~q ;
wire \always4~0_combout ;
wire \jam_reg~4_combout ;
wire \jam_reg[0]~q ;
wire \jam_reg~3_combout ;
wire \jam_reg[3]~1_combout ;
wire \jam_reg[1]~q ;
wire \jam_reg~2_combout ;
wire \jam_reg[2]~q ;
wire \jam_reg~0_combout ;
wire \jam_reg[3]~q ;
wire \tx_en_s~0_combout ;
wire \tx_en_s~1_combout ;
wire \rd_1[4]~q ;
wire \rd_2[4]~q ;
wire \rd_3[4]~q ;
wire \rd_4[4]~q ;
wire \rd_5[4]~q ;
wire \rd_6[4]~q ;
wire \always17~1_combout ;
wire \rd_7[4]~q ;
wire \rd_8[4]~q ;
wire \rd_9[4]~q ;
wire \rd_10[4]~q ;
wire \rd_11[4]~q ;
wire \rd_12[4]~q ;
wire \rd_13[6]~0_combout ;
wire \rd_13[4]~q ;
wire \always19~0_combout ;
wire \rd_14~0_combout ;
wire \rd_14[2]~1_combout ;
wire \rd_14~2_combout ;
wire \rd_1[0]~q ;
wire \rd_2[0]~q ;
wire \rd_3[0]~q ;
wire \rd_4[0]~q ;
wire \rd_5[0]~q ;
wire \rd_6[0]~q ;
wire \rd_7[0]~q ;
wire \rd_8[0]~q ;
wire \rd_9[0]~q ;
wire \rd_10[0]~q ;
wire \rd_11[0]~q ;
wire \rd_12[0]~q ;
wire \rd_13[0]~q ;
wire \rd_14~3_combout ;
wire \rd_1[5]~q ;
wire \rd_2[5]~q ;
wire \rd_3[5]~q ;
wire \rd_4[5]~q ;
wire \rd_5[5]~q ;
wire \rd_6[5]~q ;
wire \rd_7[5]~q ;
wire \rd_8[5]~q ;
wire \rd_9[5]~q ;
wire \rd_10[5]~q ;
wire \rd_11[5]~q ;
wire \rd_12[5]~q ;
wire \rd_13[5]~q ;
wire \rd_14~4_combout ;
wire \rd_1[1]~q ;
wire \rd_2[1]~q ;
wire \rd_3[1]~q ;
wire \rd_4[1]~q ;
wire \rd_5[1]~q ;
wire \rd_6[1]~q ;
wire \rd_7[1]~q ;
wire \rd_8[1]~q ;
wire \rd_9[1]~q ;
wire \rd_10[1]~q ;
wire \rd_11[1]~q ;
wire \rd_12[1]~q ;
wire \rd_13[1]~q ;
wire \rd_14~5_combout ;
wire \rd_1[6]~q ;
wire \rd_2[6]~q ;
wire \rd_3[6]~q ;
wire \rd_4[6]~q ;
wire \rd_5[6]~q ;
wire \rd_6[6]~q ;
wire \rd_7[6]~q ;
wire \rd_8[6]~q ;
wire \rd_9[6]~q ;
wire \rd_10[6]~q ;
wire \rd_11[6]~q ;
wire \rd_12[6]~q ;
wire \rd_13[6]~q ;
wire \rd_14~6_combout ;
wire \rd_1[2]~q ;
wire \rd_2[2]~q ;
wire \rd_3[2]~q ;
wire \rd_4[2]~q ;
wire \rd_5[2]~q ;
wire \rd_6[2]~q ;
wire \rd_7[2]~q ;
wire \rd_8[2]~q ;
wire \rd_9[2]~q ;
wire \rd_10[2]~q ;
wire \rd_11[2]~q ;
wire \rd_12[2]~q ;
wire \rd_13[2]~q ;
wire \rd_14~7_combout ;
wire \always19~3_wirecell_combout ;
wire \rd_1[7]~q ;
wire \rd_2[7]~q ;
wire \rd_3[7]~q ;
wire \rd_4[7]~q ;
wire \rd_5[7]~q ;
wire \rd_6[7]~q ;
wire \rd_7[7]~q ;
wire \rd_8[7]~q ;
wire \rd_9[7]~q ;
wire \rd_10[7]~q ;
wire \rd_11[7]~q ;
wire \rd_12[7]~q ;
wire \rd_13[7]~q ;
wire \rd_14~8_combout ;
wire \rd_1[3]~q ;
wire \rd_2[3]~q ;
wire \rd_3[3]~q ;
wire \rd_4[3]~q ;
wire \rd_5[3]~q ;
wire \rd_6[3]~q ;
wire \rd_7[3]~q ;
wire \rd_8[3]~q ;
wire \rd_9[3]~q ;
wire \rd_10[3]~q ;
wire \rd_11[3]~q ;
wire \rd_12[3]~q ;
wire \rd_13[3]~q ;
wire \rd_14~9_combout ;
wire \always14~0_combout ;
wire \tx_err_s[0]~q ;
wire \tx_err_s[1]~q ;
wire \tx_err_s~0_combout ;
wire \tx_err_s[2]~q ;
wire \tx_err_s[3]~q ;
wire \tx_err_s[4]~q ;
wire \tx_err_s[5]~q ;
wire \tx_err_s[6]~q ;
wire \tx_err_s[7]~q ;
wire \tx_err_s[8]~q ;
wire \tx_err_s[9]~q ;
wire \tx_err_s[10]~q ;
wire \tx_err_s[11]~q ;
wire \tx_err_s[12]~q ;
wire \tx_err_s[13]~q ;
wire \tx_err_s[14]~q ;
wire \tx_err_s[15]~q ;
wire \tx_err_s[16]~q ;
wire \tx_err_s[17]~q ;
wire \tx_err_s[18]~q ;
wire \tx_err_s[19]~q ;
wire \tx_err~0_combout ;
wire \gm_rx_crs_reg3~0_combout ;
wire \gm_rx_crs_reg3~q ;
wire \gm_rx_crs_reg4~0_combout ;
wire \gm_rx_crs_reg4~q ;
wire \frm_wait~0_combout ;
wire \tx_sav_int_reg~q ;
wire \frm_wait~1_combout ;
wire \frm_wait~2_combout ;
wire \frm_wait~3_combout ;
wire \frm_wait~q ;
wire \tx_en_s[2]~q ;
wire \tx_en_s[3]~q ;
wire \col_int~0_combout ;
wire \always9~5_combout ;
wire \always6~3_combout ;
wire \tx_stat_rden_i~q ;
wire \tx_stat_rden~0_combout ;


IoTOctopus_QSYS_altera_tse_crc328generator U_CRC(
	.txclk_ena(txclk_ena),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.sop_4(\sop[4]~q ),
	.eof_dly_5(\U_CRC|U_CTL|eof_dly[5]~q ),
	.rd_5_4(\rd_5[4]~q ),
	.rd_5_0(\rd_5[0]~q ),
	.rd_5_5(\rd_5[5]~q ),
	.rd_5_1(\rd_5[1]~q ),
	.rd_5_6(\rd_5[6]~q ),
	.rd_5_2(\rd_5[2]~q ),
	.rd_5_7(\rd_5[7]~q ),
	.rd_5_3(\rd_5[3]~q ),
	.eop_4(\eop[4]~q ),
	.reg_out_0(\U_CRC|U_GALS|reg_out[0]~_wirecell_combout ),
	.reg_out_10(\U_CRC|U_GALS|reg_out[10]~_wirecell_combout ),
	.reg_out_11(\U_CRC|U_GALS|reg_out[11]~_wirecell_combout ),
	.reg_out_12(\U_CRC|U_GALS|reg_out[12]~_wirecell_combout ),
	.reg_out_13(\U_CRC|U_GALS|reg_out[13]~_wirecell_combout ),
	.reg_out_14(\U_CRC|U_GALS|reg_out[14]~_wirecell_combout ),
	.reg_out_15(\U_CRC|U_GALS|reg_out[15]~_wirecell_combout ),
	.reg_out_16(\U_CRC|U_GALS|reg_out[16]~_wirecell_combout ),
	.reg_out_17(\U_CRC|U_GALS|reg_out[17]~_wirecell_combout ),
	.reg_out_18(\U_CRC|U_GALS|reg_out[18]~_wirecell_combout ),
	.reg_out_19(\U_CRC|U_GALS|reg_out[19]~_wirecell_combout ),
	.reg_out_1(\U_CRC|U_GALS|reg_out[1]~_wirecell_combout ),
	.reg_out_20(\U_CRC|U_GALS|reg_out[20]~_wirecell_combout ),
	.reg_out_21(\U_CRC|U_GALS|reg_out[21]~_wirecell_combout ),
	.reg_out_22(\U_CRC|U_GALS|reg_out[22]~_wirecell_combout ),
	.reg_out_23(\U_CRC|U_GALS|reg_out[23]~_wirecell_combout ),
	.reg_out_24(\U_CRC|U_GALS|reg_out[24]~_wirecell_combout ),
	.reg_out_25(\U_CRC|U_GALS|reg_out[25]~_wirecell_combout ),
	.reg_out_26(\U_CRC|U_GALS|reg_out[26]~_wirecell_combout ),
	.reg_out_27(\U_CRC|U_GALS|reg_out[27]~_wirecell_combout ),
	.reg_out_28(\U_CRC|U_GALS|reg_out[28]~_wirecell_combout ),
	.reg_out_29(\U_CRC|U_GALS|reg_out[29]~_wirecell_combout ),
	.reg_out_2(\U_CRC|U_GALS|reg_out[2]~_wirecell_combout ),
	.reg_out_30(\U_CRC|U_GALS|reg_out[30]~_wirecell_combout ),
	.reg_out_31(\U_CRC|U_GALS|reg_out[31]~_wirecell_combout ),
	.reg_out_3(\U_CRC|U_GALS|reg_out[3]~_wirecell_combout ),
	.reg_out_4(\U_CRC|U_GALS|reg_out[4]~_wirecell_combout ),
	.reg_out_5(\U_CRC|U_GALS|reg_out[5]~_wirecell_combout ),
	.reg_out_6(\U_CRC|U_GALS|reg_out[6]~_wirecell_combout ),
	.reg_out_7(\U_CRC|U_GALS|reg_out[7]~_wirecell_combout ),
	.reg_out_8(\U_CRC|U_GALS|reg_out[8]~_wirecell_combout ),
	.reg_out_9(\U_CRC|U_GALS|reg_out[9]~_wirecell_combout ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_132 U_SYNC_7(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_7|std_sync_no_cut|dreg[1]~q ),
	.gm_rx_col_reg(\gm_rx_col_reg~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_131 U_SYNC_6(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.m_rx_crs(m_rx_crs),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_9 U_SYNC_3(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_129 U_SYNC_2(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_128 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.ethernet_mode(ethernet_mode),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_134 U_SYNC_SLEEP_ENA(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_SLEEP_ENA|std_sync_no_cut|dreg[1]~q ),
	.sleep_ena(sleep_ena),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_133 U_SYNC_MAGIC_ENA(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_MAGIC_ENA|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_130 U_SYNC_4(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

dffeas gm_rx_col_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(\gm_rx_col_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\gm_rx_col_reg~q ),
	.prn(vcc));
defparam gm_rx_col_reg.is_wysiwyg = "true";
defparam gm_rx_col_reg.power_up = "low";

cyclonev_lcell_comb \gm_rx_col_reg~0 (
	.dataa(!\tx_en_s[2]~q ),
	.datab(!\gm_rx_col_reg~q ),
	.datac(!dreg_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gm_rx_col_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gm_rx_col_reg~0 .extended_lut = "off";
defparam \gm_rx_col_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \gm_rx_col_reg~0 .shared_arith = "off";

dffeas tx_ff_uflow(
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_ff_uflow~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_ff_uflow1),
	.prn(vcc));
defparam tx_ff_uflow.is_wysiwyg = "true";
defparam tx_ff_uflow.power_up = "low";

dffeas \tx_en_s[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_en_s~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(tx_en_s_1),
	.prn(vcc));
defparam \tx_en_s[1] .is_wysiwyg = "true";
defparam \tx_en_s[1] .power_up = "low";

dffeas \rd_14[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_4),
	.prn(vcc));
defparam \rd_14[4] .is_wysiwyg = "true";
defparam \rd_14[4] .power_up = "low";

dffeas \rd_14[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_0),
	.prn(vcc));
defparam \rd_14[0] .is_wysiwyg = "true";
defparam \rd_14[0] .power_up = "low";

dffeas \rd_14[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_5),
	.prn(vcc));
defparam \rd_14[5] .is_wysiwyg = "true";
defparam \rd_14[5] .power_up = "low";

dffeas \rd_14[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_1),
	.prn(vcc));
defparam \rd_14[1] .is_wysiwyg = "true";
defparam \rd_14[1] .power_up = "low";

dffeas \rd_14[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_6),
	.prn(vcc));
defparam \rd_14[6] .is_wysiwyg = "true";
defparam \rd_14[6] .power_up = "low";

dffeas \rd_14[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_2),
	.prn(vcc));
defparam \rd_14[2] .is_wysiwyg = "true";
defparam \rd_14[2] .power_up = "low";

dffeas \rd_14[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_7),
	.prn(vcc));
defparam \rd_14[7] .is_wysiwyg = "true";
defparam \rd_14[7] .power_up = "low";

dffeas \rd_14[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_14~9_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(rd_14_3),
	.prn(vcc));
defparam \rd_14[3] .is_wysiwyg = "true";
defparam \rd_14[3] .power_up = "low";

dffeas tx_err(
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_err1),
	.prn(vcc));
defparam tx_err.is_wysiwyg = "true";
defparam tx_err.power_up = "low";

cyclonev_lcell_comb \always9~1 (
	.dataa(!\frm_wait~q ),
	.datab(!\gap_wait~q ),
	.datac(!\tx_sav_int_reg~q ),
	.datad(!empty_flag),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always9),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~1 .extended_lut = "off";
defparam \always9~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \always9~1 .shared_arith = "off";

dffeas col_int(
	.clk(mac_tx_clock_connection_clk),
	.d(\col_int~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(col_int1),
	.prn(vcc));
defparam col_int.is_wysiwyg = "true";
defparam col_int.power_up = "low";

cyclonev_lcell_comb \always9~3 (
	.dataa(!q_b_9),
	.datab(!tx_data_int_7),
	.datac(!eop_sft_0),
	.datad(!\always9~0_combout ),
	.datae(!\eop_0~0_combout ),
	.dataf(!\eop_0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always91),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~3 .extended_lut = "off";
defparam \always9~3 .lut_mask = 64'hFFFFB8FFFFFFFFFF;
defparam \always9~3 .shared_arith = "off";

dffeas tx_rden_mii(
	.clk(mac_tx_clock_connection_clk),
	.d(always92),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_rden_mii1),
	.prn(vcc));
defparam tx_rden_mii.is_wysiwyg = "true";
defparam tx_rden_mii.power_up = "low";

cyclonev_lcell_comb \tx_rden_int~0 (
	.dataa(!txclk_ena),
	.datab(!dreg_1),
	.datac(!always91),
	.datad(!always9),
	.datae(!tx_rden_mii1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(tx_rden_int),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_rden_int~0 .extended_lut = "off";
defparam \tx_rden_int~0 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \tx_rden_int~0 .shared_arith = "off";

cyclonev_lcell_comb \always9~4 (
	.dataa(!\eop_0~0_combout ),
	.datab(!always9),
	.datac(!q_b_9),
	.datad(!eop_sft_0),
	.datae(!\always9~5_combout ),
	.dataf(!tx_data_int_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always92),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~4 .extended_lut = "off";
defparam \always9~4 .lut_mask = 64'hFFBBFFFFFFF3FFFF;
defparam \always9~4 .shared_arith = "off";

dffeas tx_stat_rden(
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_stat_rden~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_stat_rden1),
	.prn(vcc));
defparam tx_stat_rden.is_wysiwyg = "true";
defparam tx_stat_rden.power_up = "low";

dffeas gm_rx_col_reg2(
	.clk(mac_tx_clock_connection_clk),
	.d(\U_SYNC_7|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gm_rx_col_reg2~q ),
	.prn(vcc));
defparam gm_rx_col_reg2.is_wysiwyg = "true";
defparam gm_rx_col_reg2.power_up = "low";

cyclonev_lcell_comb \always3~0 (
	.dataa(!dreg_1),
	.datab(!\gm_rx_col_reg2~q ),
	.datac(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always3~0 .extended_lut = "off";
defparam \always3~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \always3~0 .shared_arith = "off";

cyclonev_lcell_comb \always9~0 (
	.dataa(!\frm_rd[0]~q ),
	.datab(!tx_empty),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'h7777777777777777;
defparam \always9~0 .shared_arith = "off";

cyclonev_lcell_comb \eop_0~1 (
	.dataa(!\frm_rd[2]~q ),
	.datab(!dreg_1),
	.datac(!tx_en_s_1),
	.datad(!\gm_rx_col_reg2~q ),
	.datae(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop_0~1 .extended_lut = "off";
defparam \eop_0~1 .lut_mask = 64'hFFFFFFFBFFFFFFFB;
defparam \eop_0~1 .shared_arith = "off";

cyclonev_lcell_comb \always9~2 (
	.dataa(!tx_eop_int),
	.datab(!\always9~0_combout ),
	.datac(!\eop_0~0_combout ),
	.datad(!\eop_0~1_combout ),
	.datae(!always9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~2 .extended_lut = "off";
defparam \always9~2 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \always9~2 .shared_arith = "off";

dffeas tx_rden(
	.clk(mac_tx_clock_connection_clk),
	.d(\always9~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_rden~q ),
	.prn(vcc));
defparam tx_rden.is_wysiwyg = "true";
defparam tx_rden.power_up = "low";

dffeas tx_rden_d1(
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_rden~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_rden_d1~q ),
	.prn(vcc));
defparam tx_rden_d1.is_wysiwyg = "true";
defparam tx_rden_d1.power_up = "low";

cyclonev_lcell_comb \eop_0~0 (
	.dataa(!\tx_rden~q ),
	.datab(!\tx_rden_d1~q ),
	.datac(!dreg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop_0~0 .extended_lut = "off";
defparam \eop_0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \eop_0~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_rd~0 (
	.dataa(!\always3~0_combout ),
	.datab(!tx_eop_int),
	.datac(!\always9~0_combout ),
	.datad(!\eop_0~0_combout ),
	.datae(!\eop_0~1_combout ),
	.dataf(!always9),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_rd~0 .extended_lut = "off";
defparam \frm_rd~0 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \frm_rd~0 .shared_arith = "off";

dffeas \frm_rd[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_rd~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\frm_rd[0]~q ),
	.prn(vcc));
defparam \frm_rd[0] .is_wysiwyg = "true";
defparam \frm_rd[0] .power_up = "low";

cyclonev_lcell_comb \eop_0~2 (
	.dataa(!q_b_9),
	.datab(!tx_data_int_7),
	.datac(!eop_sft_0),
	.datad(!\eop_0~0_combout ),
	.datae(!\eop_0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop_0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop_0~2 .extended_lut = "off";
defparam \eop_0~2 .lut_mask = 64'hDFFF1FFFDFFF1FFF;
defparam \eop_0~2 .shared_arith = "off";

cyclonev_lcell_comb \always6~0 (
	.dataa(!\frm_rd[0]~q ),
	.datab(!tx_empty),
	.datac(!\eop_0~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \always6~0 .shared_arith = "off";

dffeas \frm_rd[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always6~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\frm_rd[2]~q ),
	.prn(vcc));
defparam \frm_rd[2] .is_wysiwyg = "true";
defparam \frm_rd[2] .power_up = "low";

cyclonev_lcell_comb \tx_ff_uflow~0 (
	.dataa(!txclk_ena),
	.datab(!\frm_rd[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_ff_uflow~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_ff_uflow~0 .extended_lut = "off";
defparam \tx_ff_uflow~0 .lut_mask = 64'h7777777777777777;
defparam \tx_ff_uflow~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[0]~3 (
	.dataa(!txclk_ena),
	.datab(!\frm_cnt[1]~0_combout ),
	.datac(!\tx_rden~q ),
	.datad(!tx_data_int_7),
	.datae(!q_b_8),
	.dataf(!sop_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[0]~3 .extended_lut = "off";
defparam \frm_cnt[0]~3 .lut_mask = 64'hFFFFFFFFFFFFDDF5;
defparam \frm_cnt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[2]~7 (
	.dataa(!\frm_cnt[2]~q ),
	.datab(!\frm_cnt[1]~q ),
	.datac(!\frm_cnt[0]~q ),
	.datad(!\frm_cnt[4]~1_combout ),
	.datae(!\frm_cnt[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[2]~7 .extended_lut = "off";
defparam \frm_cnt[2]~7 .lut_mask = 64'hFF96FFFFFF96FFFF;
defparam \frm_cnt[2]~7 .shared_arith = "off";

dffeas \frm_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_cnt[2]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\frm_cnt[2]~q ),
	.prn(vcc));
defparam \frm_cnt[2] .is_wysiwyg = "true";
defparam \frm_cnt[2] .power_up = "low";

cyclonev_lcell_comb \frm_cnt[3]~6 (
	.dataa(!\frm_cnt[3]~q ),
	.datab(!\frm_cnt[2]~q ),
	.datac(!\frm_cnt[1]~q ),
	.datad(!\frm_cnt[0]~q ),
	.datae(!\frm_cnt[4]~1_combout ),
	.dataf(!\frm_cnt[0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[3]~6 .extended_lut = "off";
defparam \frm_cnt[3]~6 .lut_mask = 64'hFFFF6996FFFFFFFF;
defparam \frm_cnt[3]~6 .shared_arith = "off";

dffeas \frm_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_cnt[3]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\frm_cnt[3]~q ),
	.prn(vcc));
defparam \frm_cnt[3] .is_wysiwyg = "true";
defparam \frm_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\frm_cnt[3]~q ),
	.datab(!\frm_cnt[2]~q ),
	.datac(!\frm_cnt[1]~q ),
	.datad(!\frm_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[4]~5 (
	.dataa(!\frm_cnt[4]~q ),
	.datab(!\frm_cnt[4]~1_combout ),
	.datac(!\Add0~0_combout ),
	.datad(!\frm_cnt[0]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[4]~5 .extended_lut = "off";
defparam \frm_cnt[4]~5 .lut_mask = 64'hDEFFDEFFDEFFDEFF;
defparam \frm_cnt[4]~5 .shared_arith = "off";

dffeas \frm_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_cnt[4]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\frm_cnt[4]~q ),
	.prn(vcc));
defparam \frm_cnt[4] .is_wysiwyg = "true";
defparam \frm_cnt[4] .power_up = "low";

cyclonev_lcell_comb \frm_cnt[5]~4 (
	.dataa(!\frm_cnt[5]~q ),
	.datab(!\frm_cnt[4]~q ),
	.datac(!\frm_cnt[4]~1_combout ),
	.datad(!\Add0~0_combout ),
	.datae(!\frm_cnt[0]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[5]~4 .extended_lut = "off";
defparam \frm_cnt[5]~4 .lut_mask = 64'hF9F6FFFFF9F6FFFF;
defparam \frm_cnt[5]~4 .shared_arith = "off";

dffeas \frm_cnt[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_cnt[5]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\frm_cnt[5]~q ),
	.prn(vcc));
defparam \frm_cnt[5] .is_wysiwyg = "true";
defparam \frm_cnt[5] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\frm_cnt[5]~q ),
	.datab(!\frm_cnt[4]~q ),
	.datac(!\frm_cnt[3]~q ),
	.datad(!\frm_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[1]~0 (
	.dataa(!\always9~0_combout ),
	.datab(!always9),
	.datac(!\frm_cnt[1]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\frm_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[1]~0 .extended_lut = "off";
defparam \frm_cnt[1]~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \frm_cnt[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[4]~1 (
	.dataa(!txclk_ena),
	.datab(!\frm_rd[0]~q ),
	.datac(!\frm_cnt[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[4]~1 .extended_lut = "off";
defparam \frm_cnt[4]~1 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \frm_cnt[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[0]~8 (
	.dataa(!\frm_cnt[0]~q ),
	.datab(!\frm_cnt[4]~1_combout ),
	.datac(!\frm_cnt[0]~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[0]~8 .extended_lut = "off";
defparam \frm_cnt[0]~8 .lut_mask = 64'h8D8D8D8D8D8D8D8D;
defparam \frm_cnt[0]~8 .shared_arith = "off";

dffeas \frm_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_cnt[0]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\frm_cnt[0]~q ),
	.prn(vcc));
defparam \frm_cnt[0] .is_wysiwyg = "true";
defparam \frm_cnt[0] .power_up = "low";

cyclonev_lcell_comb \always6~2 (
	.dataa(!\tx_rden~q ),
	.datab(!tx_data_int_7),
	.datac(!q_b_8),
	.datad(!sop_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~2 .extended_lut = "off";
defparam \always6~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \always6~2 .shared_arith = "off";

cyclonev_lcell_comb \frm_cnt[1]~2 (
	.dataa(!\frm_cnt[1]~q ),
	.datab(!\frm_cnt[0]~q ),
	.datac(!\frm_cnt[1]~0_combout ),
	.datad(!\frm_cnt[4]~1_combout ),
	.datae(!\always6~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_cnt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_cnt[1]~2 .extended_lut = "off";
defparam \frm_cnt[1]~2 .lut_mask = 64'hF9F6FFFFF9F6FFFF;
defparam \frm_cnt[1]~2 .shared_arith = "off";

dffeas \frm_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_cnt[1]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\frm_cnt[1]~q ),
	.prn(vcc));
defparam \frm_cnt[1] .is_wysiwyg = "true";
defparam \frm_cnt[1] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\frm_cnt[5]~q ),
	.datab(!\frm_cnt[4]~q ),
	.datac(!\frm_cnt[3]~q ),
	.datad(!\frm_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \always6~1 (
	.dataa(!\frm_rd[0]~q ),
	.datab(!\eop_0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~1 .extended_lut = "off";
defparam \always6~1 .lut_mask = 64'h7777777777777777;
defparam \always6~1 .shared_arith = "off";

dffeas \frm_rd[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always6~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\frm_rd[1]~q ),
	.prn(vcc));
defparam \frm_rd[1] .is_wysiwyg = "true";
defparam \frm_rd[1] .power_up = "low";

cyclonev_lcell_comb \always7~0 (
	.dataa(!\frm_rd[1]~q ),
	.datab(!\frm_cnt[1]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\LessThan0~0_combout ),
	.datae(!\frm_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always7~0 .extended_lut = "off";
defparam \always7~0 .lut_mask = 64'hFFFFF7D5FFFFF7D5;
defparam \always7~0 .shared_arith = "off";

cyclonev_lcell_comb \pad_cnt[5]~0 (
	.dataa(!txclk_ena),
	.datab(!\always7~0_combout ),
	.datac(!\always7~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt[5]~0 .extended_lut = "off";
defparam \pad_cnt[5]~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \pad_cnt[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\pad_cnt[1]~q ),
	.datab(!\pad_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Add1~0 .shared_arith = "off";

cyclonev_lcell_comb \pad_cnt[2]~5 (
	.dataa(!col_int1),
	.datab(!\frm_cnt[2]~q ),
	.datac(!\pad_cnt[2]~q ),
	.datad(!\always7~0_combout ),
	.datae(!\pad_cnt[5]~0_combout ),
	.dataf(!\Add1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt[2]~5 .extended_lut = "off";
defparam \pad_cnt[2]~5 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \pad_cnt[2]~5 .shared_arith = "off";

dffeas \pad_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pad_cnt[2]~q ),
	.prn(vcc));
defparam \pad_cnt[2] .is_wysiwyg = "true";
defparam \pad_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\pad_cnt[2]~q ),
	.datab(!\Add1~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \pad_cnt[3]~4 (
	.dataa(!col_int1),
	.datab(!\frm_cnt[3]~q ),
	.datac(!\pad_cnt[3]~q ),
	.datad(!\always7~0_combout ),
	.datae(!\pad_cnt[5]~0_combout ),
	.dataf(!\Add1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt[3]~4 .extended_lut = "off";
defparam \pad_cnt[3]~4 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \pad_cnt[3]~4 .shared_arith = "off";

dffeas \pad_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pad_cnt[3]~q ),
	.prn(vcc));
defparam \pad_cnt[3] .is_wysiwyg = "true";
defparam \pad_cnt[3] .power_up = "low";

cyclonev_lcell_comb \pad_cnt[4]~6 (
	.dataa(!\Add1~1_combout ),
	.datab(!\pad_cnt[5]~0_combout ),
	.datac(!\frm_cnt[4]~q ),
	.datad(!\pad_cnt[4]~q ),
	.datae(!\always7~0_combout ),
	.dataf(!col_int1),
	.datag(!\pad_cnt[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt[4]~6 .extended_lut = "on";
defparam \pad_cnt[4]~6 .lut_mask = 64'h69969F6F69969F6F;
defparam \pad_cnt[4]~6 .shared_arith = "off";

dffeas \pad_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_cnt[4]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pad_cnt[4]~q ),
	.prn(vcc));
defparam \pad_cnt[4] .is_wysiwyg = "true";
defparam \pad_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Add1~2 (
	.dataa(!\pad_cnt[4]~q ),
	.datab(!\pad_cnt[3]~q ),
	.datac(!\Add1~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~2 .extended_lut = "off";
defparam \Add1~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Add1~2 .shared_arith = "off";

cyclonev_lcell_comb \pad_cnt[5]~3 (
	.dataa(!col_int1),
	.datab(!\frm_cnt[5]~q ),
	.datac(!\pad_cnt[5]~q ),
	.datad(!\always7~0_combout ),
	.datae(!\pad_cnt[5]~0_combout ),
	.dataf(!\Add1~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt[5]~3 .extended_lut = "off";
defparam \pad_cnt[5]~3 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \pad_cnt[5]~3 .shared_arith = "off";

dffeas \pad_cnt[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_cnt[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pad_cnt[5]~q ),
	.prn(vcc));
defparam \pad_cnt[5] .is_wysiwyg = "true";
defparam \pad_cnt[5] .power_up = "low";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!\pad_cnt[5]~q ),
	.datab(!\pad_cnt[4]~q ),
	.datac(!\pad_cnt[3]~q ),
	.datad(!\pad_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!\pad_cnt[5]~q ),
	.datab(!\pad_cnt[4]~q ),
	.datac(!\pad_cnt[3]~q ),
	.datad(!\pad_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \always7~1 (
	.dataa(!\pad_cnt[1]~q ),
	.datab(!\pad_cnt[0]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\Equal1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always7~1 .extended_lut = "off";
defparam \always7~1 .lut_mask = 64'h8DFF8DFF8DFF8DFF;
defparam \always7~1 .shared_arith = "off";

cyclonev_lcell_comb \pad_cnt~2 (
	.dataa(!col_int1),
	.datab(!\pad_cnt[0]~q ),
	.datac(!\frm_cnt[0]~q ),
	.datad(!\always7~0_combout ),
	.datae(!\always7~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt~2 .extended_lut = "off";
defparam \pad_cnt~2 .lut_mask = 64'hEFBFBFEFEFBFBFEF;
defparam \pad_cnt~2 .shared_arith = "off";

dffeas \pad_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_cnt~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\pad_cnt[0]~q ),
	.prn(vcc));
defparam \pad_cnt[0] .is_wysiwyg = "true";
defparam \pad_cnt[0] .power_up = "low";

cyclonev_lcell_comb \pad_cnt[1]~1 (
	.dataa(!col_int1),
	.datab(!\frm_cnt[1]~q ),
	.datac(!\pad_cnt[1]~q ),
	.datad(!\pad_cnt[0]~q ),
	.datae(!\always7~0_combout ),
	.dataf(!\pad_cnt[5]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_cnt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_cnt[1]~1 .extended_lut = "off";
defparam \pad_cnt[1]~1 .lut_mask = 64'hDFFDFDDFFDDFDFFD;
defparam \pad_cnt[1]~1 .shared_arith = "off";

dffeas \pad_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_cnt[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pad_cnt[1]~q ),
	.prn(vcc));
defparam \pad_cnt[1] .is_wysiwyg = "true";
defparam \pad_cnt[1] .power_up = "low";

cyclonev_lcell_comb \pad_wait~0 (
	.dataa(!\frm_cnt[1]~q ),
	.datab(!\Equal0~0_combout ),
	.datac(!\LessThan0~0_combout ),
	.datad(!\pad_cnt[1]~q ),
	.datae(!\pad_cnt[0]~q ),
	.dataf(!\Equal3~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pad_wait~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pad_wait~0 .extended_lut = "off";
defparam \pad_wait~0 .lut_mask = 64'hFFFFFFFFFEFDFDFE;
defparam \pad_wait~0 .shared_arith = "off";

dffeas pad_wait(
	.clk(mac_tx_clock_connection_clk),
	.d(\pad_wait~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\pad_wait~q ),
	.prn(vcc));
defparam pad_wait.is_wysiwyg = "true";
defparam pad_wait.power_up = "low";

cyclonev_lcell_comb \tx_ipg_len_int~0 (
	.dataa(!\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_ipg_len_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_ipg_len_int~0 .extended_lut = "off";
defparam \tx_ipg_len_int~0 .lut_mask = 64'hFFFFFF7DFFFFFF7D;
defparam \tx_ipg_len_int~0 .shared_arith = "off";

dffeas \tx_ipg_len_int[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_ipg_len_int~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_ipg_len_int[0]~q ),
	.prn(vcc));
defparam \tx_ipg_len_int[0] .is_wysiwyg = "true";
defparam \tx_ipg_len_int[0] .power_up = "low";

cyclonev_lcell_comb \tx_ipg_len_int~1 (
	.dataa(!\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_ipg_len_int~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_ipg_len_int~1 .extended_lut = "off";
defparam \tx_ipg_len_int~1 .lut_mask = 64'hFFBEFFFFFFBEFFFF;
defparam \tx_ipg_len_int~1 .shared_arith = "off";

dffeas \tx_ipg_len_int[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_ipg_len_int~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_ipg_len_int[1]~q ),
	.prn(vcc));
defparam \tx_ipg_len_int[1] .is_wysiwyg = "true";
defparam \tx_ipg_len_int[1] .power_up = "low";

cyclonev_lcell_comb \gap_cnt~1 (
	.dataa(!\always3~0_combout ),
	.datab(!\gap_run[4]~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\gap_cnt[0]~q ),
	.datae(!\gap_cnt[1]~q ),
	.dataf(!\tx_ipg_len_int[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gap_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gap_cnt~1 .extended_lut = "off";
defparam \gap_cnt~1 .lut_mask = 64'hBF7F7FBFFFFFFFFF;
defparam \gap_cnt~1 .shared_arith = "off";

dffeas \gap_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\gap_cnt~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_cnt[1]~q ),
	.prn(vcc));
defparam \gap_cnt[1] .is_wysiwyg = "true";
defparam \gap_cnt[1] .power_up = "low";

cyclonev_lcell_comb \tx_ipg_len_int~3 (
	.dataa(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_ipg_len_int~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_ipg_len_int~3 .extended_lut = "off";
defparam \tx_ipg_len_int~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \tx_ipg_len_int~3 .shared_arith = "off";

dffeas \tx_ipg_len_int[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_ipg_len_int~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_ipg_len_int[3]~q ),
	.prn(vcc));
defparam \tx_ipg_len_int[3] .is_wysiwyg = "true";
defparam \tx_ipg_len_int[3] .power_up = "low";

cyclonev_lcell_comb \tx_ipg_len_int~2 (
	.dataa(!\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_ipg_len_int~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_ipg_len_int~2 .extended_lut = "off";
defparam \tx_ipg_len_int~2 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \tx_ipg_len_int~2 .shared_arith = "off";

dffeas \tx_ipg_len_int[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_ipg_len_int~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_ipg_len_int[2]~q ),
	.prn(vcc));
defparam \tx_ipg_len_int[2] .is_wysiwyg = "true";
defparam \tx_ipg_len_int[2] .power_up = "low";

cyclonev_lcell_comb \Add2~1 (
	.dataa(!\gap_cnt[0]~q ),
	.datab(!\gap_cnt[1]~q ),
	.datac(!\gap_cnt[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h9696969696969696;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \gap_cnt~3 (
	.dataa(!\always3~0_combout ),
	.datab(!\gap_run[4]~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\tx_ipg_len_int[2]~q ),
	.datae(!\Add2~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gap_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gap_cnt~3 .extended_lut = "off";
defparam \gap_cnt~3 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \gap_cnt~3 .shared_arith = "off";

dffeas \gap_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\gap_cnt~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_cnt[2]~q ),
	.prn(vcc));
defparam \gap_cnt[2] .is_wysiwyg = "true";
defparam \gap_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add2~2 (
	.dataa(!\gap_cnt[0]~q ),
	.datab(!\gap_cnt[1]~q ),
	.datac(!\gap_cnt[2]~q ),
	.datad(!\gap_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~2 .extended_lut = "off";
defparam \Add2~2 .lut_mask = 64'h6996699669966996;
defparam \Add2~2 .shared_arith = "off";

cyclonev_lcell_comb \gap_cnt~4 (
	.dataa(!\always3~0_combout ),
	.datab(!\gap_run[4]~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\tx_ipg_len_int[3]~q ),
	.datae(!\Add2~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gap_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gap_cnt~4 .extended_lut = "off";
defparam \gap_cnt~4 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \gap_cnt~4 .shared_arith = "off";

dffeas \gap_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\gap_cnt~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_cnt[3]~q ),
	.prn(vcc));
defparam \gap_cnt[3] .is_wysiwyg = "true";
defparam \gap_cnt[3] .power_up = "low";

cyclonev_lcell_comb \tx_ipg_len_int~4 (
	.dataa(!\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_ipg_len_int~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_ipg_len_int~4 .extended_lut = "off";
defparam \tx_ipg_len_int~4 .lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam \tx_ipg_len_int~4 .shared_arith = "off";

dffeas \tx_ipg_len_int[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_ipg_len_int~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_ipg_len_int[4]~q ),
	.prn(vcc));
defparam \tx_ipg_len_int[4] .is_wysiwyg = "true";
defparam \tx_ipg_len_int[4] .power_up = "low";

cyclonev_lcell_comb \Add2~0 (
	.dataa(!\gap_cnt[0]~q ),
	.datab(!\gap_cnt[1]~q ),
	.datac(!\gap_cnt[2]~q ),
	.datad(!\gap_cnt[3]~q ),
	.datae(!\gap_cnt[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add2~0 .extended_lut = "off";
defparam \Add2~0 .lut_mask = 64'h9669699696696996;
defparam \Add2~0 .shared_arith = "off";

cyclonev_lcell_comb \gap_cnt~2 (
	.dataa(!\always3~0_combout ),
	.datab(!\gap_run[4]~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\tx_ipg_len_int[4]~q ),
	.datae(!\Add2~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gap_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gap_cnt~2 .extended_lut = "off";
defparam \gap_cnt~2 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \gap_cnt~2 .shared_arith = "off";

dffeas \gap_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\gap_cnt~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_cnt[4]~q ),
	.prn(vcc));
defparam \gap_cnt[4] .is_wysiwyg = "true";
defparam \gap_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!\gap_cnt[4]~q ),
	.datab(!\tx_ipg_len_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'h6666666666666666;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \always13~9 (
	.dataa(!\gap_cnt[3]~q ),
	.datab(!\gap_cnt[2]~q ),
	.datac(!\crc_fwd~q ),
	.datad(!\Equal6~0_combout ),
	.datae(!\tx_ipg_len_int[3]~q ),
	.dataf(!\tx_ipg_len_int[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~9 .extended_lut = "off";
defparam \always13~9 .lut_mask = 64'h6996966996696996;
defparam \always13~9 .shared_arith = "off";

cyclonev_lcell_comb \always13~10 (
	.dataa(!\gap_cnt[3]~q ),
	.datab(!\gap_cnt[2]~q ),
	.datac(!\crc_fwd~q ),
	.datad(!\Equal6~0_combout ),
	.datae(!\tx_ipg_len_int[3]~q ),
	.dataf(!\tx_ipg_len_int[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~10 .extended_lut = "off";
defparam \always13~10 .lut_mask = 64'h6996966996696996;
defparam \always13~10 .shared_arith = "off";

cyclonev_lcell_comb \Add4~0 (
	.dataa(!\tx_ipg_len_int[0]~q ),
	.datab(!\tx_ipg_len_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add4~0 .extended_lut = "off";
defparam \Add4~0 .lut_mask = 64'h7777777777777777;
defparam \Add4~0 .shared_arith = "off";

cyclonev_lcell_comb \always13~11 (
	.dataa(!\always13~9_combout ),
	.datab(!\always13~10_combout ),
	.datac(gnd),
	.datad(!\Add4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~11 .extended_lut = "off";
defparam \always13~11 .lut_mask = 64'h5533553355335533;
defparam \always13~11 .shared_arith = "off";

cyclonev_lcell_comb \always13~3 (
	.dataa(!\gap_cnt[0]~q ),
	.datab(!\tx_ipg_len_int[0]~q ),
	.datac(!\gap_cnt[1]~q ),
	.datad(!\tx_ipg_len_int[1]~q ),
	.datae(!\always13~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~3 .extended_lut = "off";
defparam \always13~3 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \always13~3 .shared_arith = "off";

dffeas gap_12_b(
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_12_b~q ),
	.prn(vcc));
defparam gap_12_b.is_wysiwyg = "true";
defparam gap_12_b.power_up = "low";

cyclonev_lcell_comb \always13~8 (
	.dataa(!\pad_wait~q ),
	.datab(!\gap_run[2]~q ),
	.datac(!\gap_run[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~8 .extended_lut = "off";
defparam \always13~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always13~8 .shared_arith = "off";

dffeas \gap_run[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_run[3]~q ),
	.prn(vcc));
defparam \gap_run[3] .is_wysiwyg = "true";
defparam \gap_run[3] .power_up = "low";

cyclonev_lcell_comb \always13~2 (
	.dataa(!\pad_wait~q ),
	.datab(!\gap_run[4]~q ),
	.datac(!\gap_12_b~q ),
	.datad(!\gap_run[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~2 .extended_lut = "off";
defparam \always13~2 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \always13~2 .shared_arith = "off";

dffeas \gap_run[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_run[4]~q ),
	.prn(vcc));
defparam \gap_run[4] .is_wysiwyg = "true";
defparam \gap_run[4] .power_up = "low";

cyclonev_lcell_comb \gap_cnt~0 (
	.dataa(!\always3~0_combout ),
	.datab(!\gap_run[4]~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\gap_cnt[0]~q ),
	.datae(!\tx_ipg_len_int[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gap_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gap_cnt~0 .extended_lut = "off";
defparam \gap_cnt~0 .lut_mask = 64'hBF1FFFFFBF1FFFFF;
defparam \gap_cnt~0 .shared_arith = "off";

dffeas \gap_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\gap_cnt~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_cnt[0]~q ),
	.prn(vcc));
defparam \gap_cnt[0] .is_wysiwyg = "true";
defparam \gap_cnt[0] .power_up = "low";

cyclonev_lcell_comb \always13~5 (
	.dataa(!\crc_fwd~q ),
	.datab(!\gap_cnt[2]~q ),
	.datac(!\tx_ipg_len_int[2]~q ),
	.datad(!\gap_cnt[3]~q ),
	.datae(!\tx_ipg_len_int[3]~q ),
	.dataf(!\Equal6~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~5 .extended_lut = "off";
defparam \always13~5 .lut_mask = 64'h6996966996696996;
defparam \always13~5 .shared_arith = "off";

cyclonev_lcell_comb \always13~6 (
	.dataa(!\gap_cnt[0]~q ),
	.datab(!\tx_ipg_len_int[0]~q ),
	.datac(!\gap_cnt[1]~q ),
	.datad(!\tx_ipg_len_int[1]~q ),
	.datae(!\always13~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~6 .extended_lut = "off";
defparam \always13~6 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \always13~6 .shared_arith = "off";

dffeas gap_12(
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_12~q ),
	.prn(vcc));
defparam gap_12.is_wysiwyg = "true";
defparam gap_12.power_up = "low";

cyclonev_lcell_comb \always13~7 (
	.dataa(!\gap_wait~q ),
	.datab(!\gap_run[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~7 .extended_lut = "off";
defparam \always13~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always13~7 .shared_arith = "off";

dffeas \gap_run[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_run[0]~q ),
	.prn(vcc));
defparam \gap_run[0] .is_wysiwyg = "true";
defparam \gap_run[0] .power_up = "low";

cyclonev_lcell_comb \always13~4 (
	.dataa(!\tx_rden~q ),
	.datab(!\pad_wait~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\gap_12~q ),
	.datae(!\gap_run[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~4 .extended_lut = "off";
defparam \always13~4 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \always13~4 .shared_arith = "off";

dffeas \gap_run[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_run[1]~q ),
	.prn(vcc));
defparam \gap_run[1] .is_wysiwyg = "true";
defparam \gap_run[1] .power_up = "low";

cyclonev_lcell_comb \always13~1 (
	.dataa(!\tx_rden~q ),
	.datab(!\pad_wait~q ),
	.datac(!\gap_run[1]~q ),
	.datad(!\gap_12~q ),
	.datae(!\gap_run[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~1 .extended_lut = "off";
defparam \always13~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \always13~1 .shared_arith = "off";

dffeas \gap_run[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_run[2]~q ),
	.prn(vcc));
defparam \gap_run[2] .is_wysiwyg = "true";
defparam \gap_run[2] .power_up = "low";

cyclonev_lcell_comb \always13~0 (
	.dataa(!\tx_rden~q ),
	.datab(!\gap_wait~q ),
	.datac(!\pad_wait~q ),
	.datad(!\gap_run[2]~q ),
	.datae(!\gap_run[4]~q ),
	.dataf(!\gap_12_b~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always13~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always13~0 .extended_lut = "off";
defparam \always13~0 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \always13~0 .shared_arith = "off";

dffeas gap_wait(
	.clk(mac_tx_clock_connection_clk),
	.d(\always13~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gap_wait~q ),
	.prn(vcc));
defparam gap_wait.is_wysiwyg = "true";
defparam gap_wait.power_up = "low";

cyclonev_lcell_comb \crc_fwd~0 (
	.dataa(!\tx_rden~q ),
	.datab(!\gap_wait~q ),
	.datac(!empty_flag),
	.datad(!\crc_fwd~q ),
	.datae(!tx_stat_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_fwd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_fwd~0 .extended_lut = "off";
defparam \crc_fwd~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \crc_fwd~0 .shared_arith = "off";

dffeas crc_fwd(
	.clk(mac_tx_clock_connection_clk),
	.d(\crc_fwd~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\crc_fwd~q ),
	.prn(vcc));
defparam crc_fwd.is_wysiwyg = "true";
defparam crc_fwd.power_up = "low";

cyclonev_lcell_comb \always17~0 (
	.dataa(!dreg_1),
	.datab(!tx_en_s_1),
	.datac(!\gm_rx_col_reg2~q ),
	.datad(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always17~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always17~0 .extended_lut = "off";
defparam \always17~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \always17~0 .shared_arith = "off";

cyclonev_lcell_comb \eop~13 (
	.dataa(!col_int1),
	.datab(!\pad_cnt[1]~q ),
	.datac(!\pad_cnt[0]~q ),
	.datad(!\Equal3~0_combout ),
	.datae(!\Equal1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~13 .extended_lut = "off";
defparam \eop~13 .lut_mask = 64'hBEFFFFFFBEFFFFFF;
defparam \eop~13 .shared_arith = "off";

dffeas \eop[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop_0~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[1]~q ),
	.prn(vcc));
defparam \eop[1] .is_wysiwyg = "true";
defparam \eop[1] .power_up = "low";

cyclonev_lcell_comb \eop~15 (
	.dataa(!\pad_cnt[1]~q ),
	.datab(!\pad_cnt[0]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\eop~13_combout ),
	.datae(!\eop[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~15 .extended_lut = "off";
defparam \eop~15 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \eop~15 .shared_arith = "off";

dffeas \eop[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~15_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[2]~q ),
	.prn(vcc));
defparam \eop[2] .is_wysiwyg = "true";
defparam \eop[2] .power_up = "low";

cyclonev_lcell_comb \eop~14 (
	.dataa(!\pad_cnt[1]~q ),
	.datab(!\pad_cnt[0]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\eop[2]~q ),
	.datae(!\eop~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~14 .extended_lut = "off";
defparam \eop~14 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \eop~14 .shared_arith = "off";

dffeas \eop[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~14_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[3]~q ),
	.prn(vcc));
defparam \eop[3] .is_wysiwyg = "true";
defparam \eop[3] .power_up = "low";

dffeas \eop[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\eop[4]~q ),
	.prn(vcc));
defparam \eop[4] .is_wysiwyg = "true";
defparam \eop[4] .power_up = "low";

cyclonev_lcell_comb \eop~12 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~12 .extended_lut = "off";
defparam \eop~12 .lut_mask = 64'h7777777777777777;
defparam \eop~12 .shared_arith = "off";

dffeas \eop[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~12_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[5]~q ),
	.prn(vcc));
defparam \eop[5] .is_wysiwyg = "true";
defparam \eop[5] .power_up = "low";

cyclonev_lcell_comb \eop~11 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~11 .extended_lut = "off";
defparam \eop~11 .lut_mask = 64'h7777777777777777;
defparam \eop~11 .shared_arith = "off";

dffeas \eop[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~11_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[6]~q ),
	.prn(vcc));
defparam \eop[6] .is_wysiwyg = "true";
defparam \eop[6] .power_up = "low";

cyclonev_lcell_comb \eop~10 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~10 .extended_lut = "off";
defparam \eop~10 .lut_mask = 64'h7777777777777777;
defparam \eop~10 .shared_arith = "off";

dffeas \eop[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~10_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[7]~q ),
	.prn(vcc));
defparam \eop[7] .is_wysiwyg = "true";
defparam \eop[7] .power_up = "low";

cyclonev_lcell_comb \eop~9 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~9 .extended_lut = "off";
defparam \eop~9 .lut_mask = 64'h7777777777777777;
defparam \eop~9 .shared_arith = "off";

dffeas \eop[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~9_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[8]~q ),
	.prn(vcc));
defparam \eop[8] .is_wysiwyg = "true";
defparam \eop[8] .power_up = "low";

cyclonev_lcell_comb \eop~8 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~8 .extended_lut = "off";
defparam \eop~8 .lut_mask = 64'h7777777777777777;
defparam \eop~8 .shared_arith = "off";

dffeas \eop[9] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[9]~q ),
	.prn(vcc));
defparam \eop[9] .is_wysiwyg = "true";
defparam \eop[9] .power_up = "low";

cyclonev_lcell_comb \eop~6 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~6 .extended_lut = "off";
defparam \eop~6 .lut_mask = 64'h7777777777777777;
defparam \eop~6 .shared_arith = "off";

dffeas \eop[10] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[10]~q ),
	.prn(vcc));
defparam \eop[10] .is_wysiwyg = "true";
defparam \eop[10] .power_up = "low";

cyclonev_lcell_comb \eop~4 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~4 .extended_lut = "off";
defparam \eop~4 .lut_mask = 64'h7777777777777777;
defparam \eop~4 .shared_arith = "off";

dffeas \eop[11] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[11]~q ),
	.prn(vcc));
defparam \eop[11] .is_wysiwyg = "true";
defparam \eop[11] .power_up = "low";

cyclonev_lcell_comb \eop~2 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~2 .extended_lut = "off";
defparam \eop~2 .lut_mask = 64'h7777777777777777;
defparam \eop~2 .shared_arith = "off";

dffeas \eop[12] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[12]~q ),
	.prn(vcc));
defparam \eop[12] .is_wysiwyg = "true";
defparam \eop[12] .power_up = "low";

cyclonev_lcell_comb \eop~0 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~0 .extended_lut = "off";
defparam \eop~0 .lut_mask = 64'h7777777777777777;
defparam \eop~0 .shared_arith = "off";

dffeas \eop[13] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[13]~q ),
	.prn(vcc));
defparam \eop[13] .is_wysiwyg = "true";
defparam \eop[13] .power_up = "low";

cyclonev_lcell_comb \eop~7 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~7 .extended_lut = "off";
defparam \eop~7 .lut_mask = 64'h7777777777777777;
defparam \eop~7 .shared_arith = "off";

dffeas \eop[14] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[14]~q ),
	.prn(vcc));
defparam \eop[14] .is_wysiwyg = "true";
defparam \eop[14] .power_up = "low";

cyclonev_lcell_comb \eop~5 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~5 .extended_lut = "off";
defparam \eop~5 .lut_mask = 64'h7777777777777777;
defparam \eop~5 .shared_arith = "off";

dffeas \eop[15] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[15]~q ),
	.prn(vcc));
defparam \eop[15] .is_wysiwyg = "true";
defparam \eop[15] .power_up = "low";

cyclonev_lcell_comb \eop~3 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~3 .extended_lut = "off";
defparam \eop~3 .lut_mask = 64'h7777777777777777;
defparam \eop~3 .shared_arith = "off";

dffeas \eop[16] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[16]~q ),
	.prn(vcc));
defparam \eop[16] .is_wysiwyg = "true";
defparam \eop[16] .power_up = "low";

cyclonev_lcell_comb \eop~1 (
	.dataa(!\always17~0_combout ),
	.datab(!\eop[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop~1 .extended_lut = "off";
defparam \eop~1 .lut_mask = 64'h7777777777777777;
defparam \eop~1 .shared_arith = "off";

dffeas \eop[17] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\eop[17]~q ),
	.prn(vcc));
defparam \eop[17] .is_wysiwyg = "true";
defparam \eop[17] .power_up = "low";

cyclonev_lcell_comb \tx_en_s~2 (
	.dataa(!\tx_en_s[0]~q ),
	.datab(!\crc_fwd~q ),
	.datac(!\eop[13]~q ),
	.datad(!\eop[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_en_s~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_en_s~2 .extended_lut = "off";
defparam \tx_en_s~2 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \tx_en_s~2 .shared_arith = "off";

cyclonev_lcell_comb \sop~0 (
	.dataa(!\sop[4]~q ),
	.datab(!\sop[3]~q ),
	.datac(!\always6~2_combout ),
	.datad(!\sop[2]~q ),
	.datae(!\sop[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop~0 .extended_lut = "off";
defparam \sop~0 .lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam \sop~0 .shared_arith = "off";

dffeas \sop[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\sop~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\sop[1]~q ),
	.prn(vcc));
defparam \sop[1] .is_wysiwyg = "true";
defparam \sop[1] .power_up = "low";

dffeas \sop[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\sop[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\sop[2]~q ),
	.prn(vcc));
defparam \sop[2] .is_wysiwyg = "true";
defparam \sop[2] .power_up = "low";

dffeas \sop[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\sop[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\sop[3]~q ),
	.prn(vcc));
defparam \sop[3] .is_wysiwyg = "true";
defparam \sop[3] .power_up = "low";

dffeas \sop[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\sop[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sop[4]~q ),
	.prn(vcc));
defparam \sop[4] .is_wysiwyg = "true";
defparam \sop[4] .power_up = "low";

dffeas \tx_en_s[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_en_s~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\sop[4]~q ),
	.ena(txclk_ena),
	.q(\tx_en_s[0]~q ),
	.prn(vcc));
defparam \tx_en_s[0] .is_wysiwyg = "true";
defparam \tx_en_s[0] .power_up = "low";

cyclonev_lcell_comb \preamb_cnt~2 (
	.dataa(!\preamb_wait~q ),
	.datab(!\preamb_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\preamb_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \preamb_cnt~2 .extended_lut = "off";
defparam \preamb_cnt~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \preamb_cnt~2 .shared_arith = "off";

dffeas \preamb_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\preamb_cnt~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_cnt[0]~q ),
	.prn(vcc));
defparam \preamb_cnt[0] .is_wysiwyg = "true";
defparam \preamb_cnt[0] .power_up = "low";

cyclonev_lcell_comb \preamb_cnt~1 (
	.dataa(!\preamb_wait~q ),
	.datab(!\preamb_cnt[1]~q ),
	.datac(!\preamb_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\preamb_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \preamb_cnt~1 .extended_lut = "off";
defparam \preamb_cnt~1 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \preamb_cnt~1 .shared_arith = "off";

dffeas \preamb_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\preamb_cnt~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_cnt[1]~q ),
	.prn(vcc));
defparam \preamb_cnt[1] .is_wysiwyg = "true";
defparam \preamb_cnt[1] .power_up = "low";

cyclonev_lcell_comb \preamb_cnt~0 (
	.dataa(!\preamb_wait~q ),
	.datab(!\preamb_cnt[2]~q ),
	.datac(!\preamb_cnt[1]~q ),
	.datad(!\preamb_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\preamb_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \preamb_cnt~0 .extended_lut = "off";
defparam \preamb_cnt~0 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \preamb_cnt~0 .shared_arith = "off";

dffeas \preamb_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\preamb_cnt~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_cnt[2]~q ),
	.prn(vcc));
defparam \preamb_cnt[2] .is_wysiwyg = "true";
defparam \preamb_cnt[2] .power_up = "low";

cyclonev_lcell_comb \always19~3 (
	.dataa(!\preamb_wait~q ),
	.datab(!\sop[4]~q ),
	.datac(!\preamb_run[0]~q ),
	.datad(!\preamb_cnt[2]~q ),
	.datae(!\preamb_cnt[1]~q ),
	.dataf(!\preamb_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always19~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always19~3 .extended_lut = "off";
defparam \always19~3 .lut_mask = 64'hFFFFFFBFFFFFFFFF;
defparam \always19~3 .shared_arith = "off";

dffeas \preamb_run[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always19~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_run[0]~q ),
	.prn(vcc));
defparam \preamb_run[0] .is_wysiwyg = "true";
defparam \preamb_run[0] .power_up = "low";

cyclonev_lcell_comb \always19~4 (
	.dataa(!\preamb_run[0]~q ),
	.datab(!\preamb_cnt[2]~q ),
	.datac(!\preamb_cnt[1]~q ),
	.datad(!\preamb_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always19~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always19~4 .extended_lut = "off";
defparam \always19~4 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \always19~4 .shared_arith = "off";

dffeas \preamb_run[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always19~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_run[1]~q ),
	.prn(vcc));
defparam \preamb_run[1] .is_wysiwyg = "true";
defparam \preamb_run[1] .power_up = "low";

cyclonev_lcell_comb \always19~2 (
	.dataa(!\preamb_run[2]~q ),
	.datab(!\crc_fwd~q ),
	.datac(!\eop[13]~q ),
	.datad(!\eop[17]~q ),
	.datae(!\preamb_run[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always19~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always19~2 .extended_lut = "off";
defparam \always19~2 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \always19~2 .shared_arith = "off";

dffeas \preamb_run[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always19~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_run[2]~q ),
	.prn(vcc));
defparam \preamb_run[2] .is_wysiwyg = "true";
defparam \preamb_run[2] .power_up = "low";

cyclonev_lcell_comb \always19~1 (
	.dataa(!\preamb_wait~q ),
	.datab(!\preamb_run[2]~q ),
	.datac(!\crc_fwd~q ),
	.datad(!\eop[13]~q ),
	.datae(!\eop[17]~q ),
	.dataf(!\sop[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always19~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always19~1 .extended_lut = "off";
defparam \always19~1 .lut_mask = 64'hBFFFFFFFB3FFFFFF;
defparam \always19~1 .shared_arith = "off";

cyclonev_lcell_comb \preamb_wait~0 (
	.dataa(!\always19~1_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\preamb_wait~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \preamb_wait~0 .extended_lut = "off";
defparam \preamb_wait~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \preamb_wait~0 .shared_arith = "off";

dffeas preamb_wait(
	.clk(mac_tx_clock_connection_clk),
	.d(\preamb_wait~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\preamb_wait~q ),
	.prn(vcc));
defparam preamb_wait.is_wysiwyg = "true";
defparam preamb_wait.power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!\gm_rx_col_reg2~q ),
	.datab(!\tx_en_s[0]~q ),
	.datac(!\U_SYNC_7|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \always4~0 .shared_arith = "off";

cyclonev_lcell_comb \jam_reg~4 (
	.dataa(!\jam_reg[0]~q ),
	.datab(!\preamb_wait~q ),
	.datac(!\preamb_run[2]~q ),
	.datad(!\always4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jam_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jam_reg~4 .extended_lut = "off";
defparam \jam_reg~4 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \jam_reg~4 .shared_arith = "off";

dffeas \jam_reg[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\jam_reg~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\jam_reg[0]~q ),
	.prn(vcc));
defparam \jam_reg[0] .is_wysiwyg = "true";
defparam \jam_reg[0] .power_up = "low";

cyclonev_lcell_comb \jam_reg~3 (
	.dataa(!\jam_reg[0]~q ),
	.datab(!\always4~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jam_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jam_reg~3 .extended_lut = "off";
defparam \jam_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \jam_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \jam_reg[3]~1 (
	.dataa(!txclk_ena),
	.datab(!\preamb_wait~q ),
	.datac(!\preamb_run[2]~q ),
	.datad(!\always4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jam_reg[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jam_reg[3]~1 .extended_lut = "off";
defparam \jam_reg[3]~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \jam_reg[3]~1 .shared_arith = "off";

dffeas \jam_reg[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\jam_reg~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jam_reg[3]~1_combout ),
	.q(\jam_reg[1]~q ),
	.prn(vcc));
defparam \jam_reg[1] .is_wysiwyg = "true";
defparam \jam_reg[1] .power_up = "low";

cyclonev_lcell_comb \jam_reg~2 (
	.dataa(!\jam_reg[1]~q ),
	.datab(!\always4~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jam_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jam_reg~2 .extended_lut = "off";
defparam \jam_reg~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \jam_reg~2 .shared_arith = "off";

dffeas \jam_reg[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\jam_reg~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jam_reg[3]~1_combout ),
	.q(\jam_reg[2]~q ),
	.prn(vcc));
defparam \jam_reg[2] .is_wysiwyg = "true";
defparam \jam_reg[2] .power_up = "low";

cyclonev_lcell_comb \jam_reg~0 (
	.dataa(!\jam_reg[2]~q ),
	.datab(!\always4~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jam_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jam_reg~0 .extended_lut = "off";
defparam \jam_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \jam_reg~0 .shared_arith = "off";

dffeas \jam_reg[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\jam_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jam_reg[3]~1_combout ),
	.q(\jam_reg[3]~q ),
	.prn(vcc));
defparam \jam_reg[3] .is_wysiwyg = "true";
defparam \jam_reg[3] .power_up = "low";

cyclonev_lcell_comb \tx_en_s~0 (
	.dataa(!\jam_reg[3]~q ),
	.datab(!\jam_reg[2]~q ),
	.datac(!\jam_reg[1]~q ),
	.datad(!\jam_reg[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_en_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_en_s~0 .extended_lut = "off";
defparam \tx_en_s~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \tx_en_s~0 .shared_arith = "off";

cyclonev_lcell_comb \tx_en_s~1 (
	.dataa(!dreg_1),
	.datab(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datac(!\tx_en_s[0]~q ),
	.datad(!\tx_en_s~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_en_s~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_en_s~1 .extended_lut = "off";
defparam \tx_en_s~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \tx_en_s~1 .shared_arith = "off";

dffeas \rd_1[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_4),
	.asdata(dout_reg_sft_28),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[4]~q ),
	.prn(vcc));
defparam \rd_1[4] .is_wysiwyg = "true";
defparam \rd_1[4] .power_up = "low";

dffeas \rd_2[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[4]~q ),
	.prn(vcc));
defparam \rd_2[4] .is_wysiwyg = "true";
defparam \rd_2[4] .power_up = "low";

dffeas \rd_3[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[4]~q ),
	.prn(vcc));
defparam \rd_3[4] .is_wysiwyg = "true";
defparam \rd_3[4] .power_up = "low";

dffeas \rd_4[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[4]~q ),
	.prn(vcc));
defparam \rd_4[4] .is_wysiwyg = "true";
defparam \rd_4[4] .power_up = "low";

dffeas \rd_5[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[4]~q ),
	.prn(vcc));
defparam \rd_5[4] .is_wysiwyg = "true";
defparam \rd_5[4] .power_up = "low";

dffeas \rd_6[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[4]~q ),
	.prn(vcc));
defparam \rd_6[4] .is_wysiwyg = "true";
defparam \rd_6[4] .power_up = "low";

cyclonev_lcell_comb \always17~1 (
	.dataa(!\crc_fwd~q ),
	.datab(!\U_CRC|U_CTL|eof_dly[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always17~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always17~1 .extended_lut = "off";
defparam \always17~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always17~1 .shared_arith = "off";

dffeas \rd_7[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[28]~_wirecell_combout ),
	.asdata(\rd_6[4]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[4]~q ),
	.prn(vcc));
defparam \rd_7[4] .is_wysiwyg = "true";
defparam \rd_7[4] .power_up = "low";

dffeas \rd_8[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[20]~_wirecell_combout ),
	.asdata(\rd_7[4]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[4]~q ),
	.prn(vcc));
defparam \rd_8[4] .is_wysiwyg = "true";
defparam \rd_8[4] .power_up = "low";

dffeas \rd_9[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[12]~_wirecell_combout ),
	.asdata(\rd_8[4]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[4]~q ),
	.prn(vcc));
defparam \rd_9[4] .is_wysiwyg = "true";
defparam \rd_9[4] .power_up = "low";

dffeas \rd_10[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[4]~_wirecell_combout ),
	.asdata(\rd_9[4]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[4]~q ),
	.prn(vcc));
defparam \rd_10[4] .is_wysiwyg = "true";
defparam \rd_10[4] .power_up = "low";

dffeas \rd_11[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[4]~q ),
	.prn(vcc));
defparam \rd_11[4] .is_wysiwyg = "true";
defparam \rd_11[4] .power_up = "low";

dffeas \rd_12[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[4]~q ),
	.prn(vcc));
defparam \rd_12[4] .is_wysiwyg = "true";
defparam \rd_12[4] .power_up = "low";

cyclonev_lcell_comb \rd_13[6]~0 (
	.dataa(!\preamb_wait~q ),
	.datab(!\sop[4]~q ),
	.datac(!\preamb_run[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_13[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_13[6]~0 .extended_lut = "off";
defparam \rd_13[6]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \rd_13[6]~0 .shared_arith = "off";

dffeas \rd_13[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(vcc),
	.asdata(\rd_12[4]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[4]~q ),
	.prn(vcc));
defparam \rd_13[4] .is_wysiwyg = "true";
defparam \rd_13[4] .power_up = "low";

cyclonev_lcell_comb \always19~0 (
	.dataa(!\jam_reg[0]~q ),
	.datab(!\preamb_wait~q ),
	.datac(!\preamb_run[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always19~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always19~0 .extended_lut = "off";
defparam \always19~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \always19~0 .shared_arith = "off";

cyclonev_lcell_comb \rd_14~0 (
	.dataa(!\jam_reg[1]~q ),
	.datab(!\always19~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~0 .extended_lut = "off";
defparam \rd_14~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \rd_14~0 .shared_arith = "off";

cyclonev_lcell_comb \rd_14[2]~1 (
	.dataa(!dreg_1),
	.datab(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datac(!\jam_reg[3]~q ),
	.datad(!\jam_reg[2]~q ),
	.datae(!\rd_14~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14[2]~1 .extended_lut = "off";
defparam \rd_14[2]~1 .lut_mask = 64'hFFFFBFFFFFFFBFFF;
defparam \rd_14[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \rd_14~2 (
	.dataa(!\jam_reg[1]~q ),
	.datab(!\rd_13[4]~q ),
	.datac(!\always19~0_combout ),
	.datad(!\rd_14[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~2 .extended_lut = "off";
defparam \rd_14~2 .lut_mask = 64'hF377F377F377F377;
defparam \rd_14~2 .shared_arith = "off";

dffeas \rd_1[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_0),
	.asdata(dout_reg_sft_24),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[0]~q ),
	.prn(vcc));
defparam \rd_1[0] .is_wysiwyg = "true";
defparam \rd_1[0] .power_up = "low";

dffeas \rd_2[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[0]~q ),
	.prn(vcc));
defparam \rd_2[0] .is_wysiwyg = "true";
defparam \rd_2[0] .power_up = "low";

dffeas \rd_3[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[0]~q ),
	.prn(vcc));
defparam \rd_3[0] .is_wysiwyg = "true";
defparam \rd_3[0] .power_up = "low";

dffeas \rd_4[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[0]~q ),
	.prn(vcc));
defparam \rd_4[0] .is_wysiwyg = "true";
defparam \rd_4[0] .power_up = "low";

dffeas \rd_5[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[0]~q ),
	.prn(vcc));
defparam \rd_5[0] .is_wysiwyg = "true";
defparam \rd_5[0] .power_up = "low";

dffeas \rd_6[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[0]~q ),
	.prn(vcc));
defparam \rd_6[0] .is_wysiwyg = "true";
defparam \rd_6[0] .power_up = "low";

dffeas \rd_7[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[24]~_wirecell_combout ),
	.asdata(\rd_6[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[0]~q ),
	.prn(vcc));
defparam \rd_7[0] .is_wysiwyg = "true";
defparam \rd_7[0] .power_up = "low";

dffeas \rd_8[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[16]~_wirecell_combout ),
	.asdata(\rd_7[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[0]~q ),
	.prn(vcc));
defparam \rd_8[0] .is_wysiwyg = "true";
defparam \rd_8[0] .power_up = "low";

dffeas \rd_9[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[8]~_wirecell_combout ),
	.asdata(\rd_8[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[0]~q ),
	.prn(vcc));
defparam \rd_9[0] .is_wysiwyg = "true";
defparam \rd_9[0] .power_up = "low";

dffeas \rd_10[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[0]~_wirecell_combout ),
	.asdata(\rd_9[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[0]~q ),
	.prn(vcc));
defparam \rd_10[0] .is_wysiwyg = "true";
defparam \rd_10[0] .power_up = "low";

dffeas \rd_11[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[0]~q ),
	.prn(vcc));
defparam \rd_11[0] .is_wysiwyg = "true";
defparam \rd_11[0] .power_up = "low";

dffeas \rd_12[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[0]~q ),
	.prn(vcc));
defparam \rd_12[0] .is_wysiwyg = "true";
defparam \rd_12[0] .power_up = "low";

dffeas \rd_13[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(vcc),
	.asdata(\rd_12[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[0]~q ),
	.prn(vcc));
defparam \rd_13[0] .is_wysiwyg = "true";
defparam \rd_13[0] .power_up = "low";

cyclonev_lcell_comb \rd_14~3 (
	.dataa(!\jam_reg[2]~q ),
	.datab(!\rd_14~0_combout ),
	.datac(!\rd_14[2]~1_combout ),
	.datad(!\rd_13[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~3 .extended_lut = "off";
defparam \rd_14~3 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \rd_14~3 .shared_arith = "off";

dffeas \rd_1[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_5),
	.asdata(dout_reg_sft_29),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[5]~q ),
	.prn(vcc));
defparam \rd_1[5] .is_wysiwyg = "true";
defparam \rd_1[5] .power_up = "low";

dffeas \rd_2[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[5]~q ),
	.prn(vcc));
defparam \rd_2[5] .is_wysiwyg = "true";
defparam \rd_2[5] .power_up = "low";

dffeas \rd_3[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[5]~q ),
	.prn(vcc));
defparam \rd_3[5] .is_wysiwyg = "true";
defparam \rd_3[5] .power_up = "low";

dffeas \rd_4[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[5]~q ),
	.prn(vcc));
defparam \rd_4[5] .is_wysiwyg = "true";
defparam \rd_4[5] .power_up = "low";

dffeas \rd_5[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[5]~q ),
	.prn(vcc));
defparam \rd_5[5] .is_wysiwyg = "true";
defparam \rd_5[5] .power_up = "low";

dffeas \rd_6[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[5]~q ),
	.prn(vcc));
defparam \rd_6[5] .is_wysiwyg = "true";
defparam \rd_6[5] .power_up = "low";

dffeas \rd_7[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[29]~_wirecell_combout ),
	.asdata(\rd_6[5]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[5]~q ),
	.prn(vcc));
defparam \rd_7[5] .is_wysiwyg = "true";
defparam \rd_7[5] .power_up = "low";

dffeas \rd_8[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[21]~_wirecell_combout ),
	.asdata(\rd_7[5]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[5]~q ),
	.prn(vcc));
defparam \rd_8[5] .is_wysiwyg = "true";
defparam \rd_8[5] .power_up = "low";

dffeas \rd_9[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[13]~_wirecell_combout ),
	.asdata(\rd_8[5]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[5]~q ),
	.prn(vcc));
defparam \rd_9[5] .is_wysiwyg = "true";
defparam \rd_9[5] .power_up = "low";

dffeas \rd_10[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[5]~_wirecell_combout ),
	.asdata(\rd_9[5]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[5]~q ),
	.prn(vcc));
defparam \rd_10[5] .is_wysiwyg = "true";
defparam \rd_10[5] .power_up = "low";

dffeas \rd_11[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[5]~q ),
	.prn(vcc));
defparam \rd_11[5] .is_wysiwyg = "true";
defparam \rd_11[5] .power_up = "low";

dffeas \rd_12[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[5]~q ),
	.prn(vcc));
defparam \rd_12[5] .is_wysiwyg = "true";
defparam \rd_12[5] .power_up = "low";

dffeas \rd_13[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rd_12[5]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[5]~q ),
	.prn(vcc));
defparam \rd_13[5] .is_wysiwyg = "true";
defparam \rd_13[5] .power_up = "low";

cyclonev_lcell_comb \rd_14~4 (
	.dataa(!\jam_reg[2]~q ),
	.datab(!\rd_14~0_combout ),
	.datac(!\rd_14[2]~1_combout ),
	.datad(!\rd_13[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~4 .extended_lut = "off";
defparam \rd_14~4 .lut_mask = 64'hACFFACFFACFFACFF;
defparam \rd_14~4 .shared_arith = "off";

dffeas \rd_1[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_1),
	.asdata(dout_reg_sft_25),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[1]~q ),
	.prn(vcc));
defparam \rd_1[1] .is_wysiwyg = "true";
defparam \rd_1[1] .power_up = "low";

dffeas \rd_2[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[1]~q ),
	.prn(vcc));
defparam \rd_2[1] .is_wysiwyg = "true";
defparam \rd_2[1] .power_up = "low";

dffeas \rd_3[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[1]~q ),
	.prn(vcc));
defparam \rd_3[1] .is_wysiwyg = "true";
defparam \rd_3[1] .power_up = "low";

dffeas \rd_4[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[1]~q ),
	.prn(vcc));
defparam \rd_4[1] .is_wysiwyg = "true";
defparam \rd_4[1] .power_up = "low";

dffeas \rd_5[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[1]~q ),
	.prn(vcc));
defparam \rd_5[1] .is_wysiwyg = "true";
defparam \rd_5[1] .power_up = "low";

dffeas \rd_6[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[1]~q ),
	.prn(vcc));
defparam \rd_6[1] .is_wysiwyg = "true";
defparam \rd_6[1] .power_up = "low";

dffeas \rd_7[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[25]~_wirecell_combout ),
	.asdata(\rd_6[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[1]~q ),
	.prn(vcc));
defparam \rd_7[1] .is_wysiwyg = "true";
defparam \rd_7[1] .power_up = "low";

dffeas \rd_8[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[17]~_wirecell_combout ),
	.asdata(\rd_7[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[1]~q ),
	.prn(vcc));
defparam \rd_8[1] .is_wysiwyg = "true";
defparam \rd_8[1] .power_up = "low";

dffeas \rd_9[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[9]~_wirecell_combout ),
	.asdata(\rd_8[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[1]~q ),
	.prn(vcc));
defparam \rd_9[1] .is_wysiwyg = "true";
defparam \rd_9[1] .power_up = "low";

dffeas \rd_10[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[1]~_wirecell_combout ),
	.asdata(\rd_9[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[1]~q ),
	.prn(vcc));
defparam \rd_10[1] .is_wysiwyg = "true";
defparam \rd_10[1] .power_up = "low";

dffeas \rd_11[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[1]~q ),
	.prn(vcc));
defparam \rd_11[1] .is_wysiwyg = "true";
defparam \rd_11[1] .power_up = "low";

dffeas \rd_12[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[1]~q ),
	.prn(vcc));
defparam \rd_12[1] .is_wysiwyg = "true";
defparam \rd_12[1] .power_up = "low";

dffeas \rd_13[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rd_12[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[1]~q ),
	.prn(vcc));
defparam \rd_13[1] .is_wysiwyg = "true";
defparam \rd_13[1] .power_up = "low";

cyclonev_lcell_comb \rd_14~5 (
	.dataa(!\rd_14~0_combout ),
	.datab(!\rd_14[2]~1_combout ),
	.datac(!\rd_13[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~5 .extended_lut = "off";
defparam \rd_14~5 .lut_mask = 64'h8B8B8B8B8B8B8B8B;
defparam \rd_14~5 .shared_arith = "off";

dffeas \rd_1[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_6),
	.asdata(dout_reg_sft_30),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[6]~q ),
	.prn(vcc));
defparam \rd_1[6] .is_wysiwyg = "true";
defparam \rd_1[6] .power_up = "low";

dffeas \rd_2[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[6]~q ),
	.prn(vcc));
defparam \rd_2[6] .is_wysiwyg = "true";
defparam \rd_2[6] .power_up = "low";

dffeas \rd_3[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[6]~q ),
	.prn(vcc));
defparam \rd_3[6] .is_wysiwyg = "true";
defparam \rd_3[6] .power_up = "low";

dffeas \rd_4[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[6]~q ),
	.prn(vcc));
defparam \rd_4[6] .is_wysiwyg = "true";
defparam \rd_4[6] .power_up = "low";

dffeas \rd_5[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[6]~q ),
	.prn(vcc));
defparam \rd_5[6] .is_wysiwyg = "true";
defparam \rd_5[6] .power_up = "low";

dffeas \rd_6[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[6]~q ),
	.prn(vcc));
defparam \rd_6[6] .is_wysiwyg = "true";
defparam \rd_6[6] .power_up = "low";

dffeas \rd_7[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[30]~_wirecell_combout ),
	.asdata(\rd_6[6]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[6]~q ),
	.prn(vcc));
defparam \rd_7[6] .is_wysiwyg = "true";
defparam \rd_7[6] .power_up = "low";

dffeas \rd_8[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[22]~_wirecell_combout ),
	.asdata(\rd_7[6]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[6]~q ),
	.prn(vcc));
defparam \rd_8[6] .is_wysiwyg = "true";
defparam \rd_8[6] .power_up = "low";

dffeas \rd_9[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[14]~_wirecell_combout ),
	.asdata(\rd_8[6]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[6]~q ),
	.prn(vcc));
defparam \rd_9[6] .is_wysiwyg = "true";
defparam \rd_9[6] .power_up = "low";

dffeas \rd_10[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[6]~_wirecell_combout ),
	.asdata(\rd_9[6]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[6]~q ),
	.prn(vcc));
defparam \rd_10[6] .is_wysiwyg = "true";
defparam \rd_10[6] .power_up = "low";

dffeas \rd_11[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[6]~q ),
	.prn(vcc));
defparam \rd_11[6] .is_wysiwyg = "true";
defparam \rd_11[6] .power_up = "low";

dffeas \rd_12[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[6]~q ),
	.prn(vcc));
defparam \rd_12[6] .is_wysiwyg = "true";
defparam \rd_12[6] .power_up = "low";

dffeas \rd_13[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(vcc),
	.asdata(\rd_12[6]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[6]~q ),
	.prn(vcc));
defparam \rd_13[6] .is_wysiwyg = "true";
defparam \rd_13[6] .power_up = "low";

cyclonev_lcell_comb \rd_14~6 (
	.dataa(!\jam_reg[2]~q ),
	.datab(!\rd_14~0_combout ),
	.datac(!\rd_14[2]~1_combout ),
	.datad(!\rd_13[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~6 .extended_lut = "off";
defparam \rd_14~6 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \rd_14~6 .shared_arith = "off";

dffeas \rd_1[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_2),
	.asdata(dout_reg_sft_26),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[2]~q ),
	.prn(vcc));
defparam \rd_1[2] .is_wysiwyg = "true";
defparam \rd_1[2] .power_up = "low";

dffeas \rd_2[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[2]~q ),
	.prn(vcc));
defparam \rd_2[2] .is_wysiwyg = "true";
defparam \rd_2[2] .power_up = "low";

dffeas \rd_3[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[2]~q ),
	.prn(vcc));
defparam \rd_3[2] .is_wysiwyg = "true";
defparam \rd_3[2] .power_up = "low";

dffeas \rd_4[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[2]~q ),
	.prn(vcc));
defparam \rd_4[2] .is_wysiwyg = "true";
defparam \rd_4[2] .power_up = "low";

dffeas \rd_5[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[2]~q ),
	.prn(vcc));
defparam \rd_5[2] .is_wysiwyg = "true";
defparam \rd_5[2] .power_up = "low";

dffeas \rd_6[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[2]~q ),
	.prn(vcc));
defparam \rd_6[2] .is_wysiwyg = "true";
defparam \rd_6[2] .power_up = "low";

dffeas \rd_7[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[26]~_wirecell_combout ),
	.asdata(\rd_6[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[2]~q ),
	.prn(vcc));
defparam \rd_7[2] .is_wysiwyg = "true";
defparam \rd_7[2] .power_up = "low";

dffeas \rd_8[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[18]~_wirecell_combout ),
	.asdata(\rd_7[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[2]~q ),
	.prn(vcc));
defparam \rd_8[2] .is_wysiwyg = "true";
defparam \rd_8[2] .power_up = "low";

dffeas \rd_9[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[10]~_wirecell_combout ),
	.asdata(\rd_8[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[2]~q ),
	.prn(vcc));
defparam \rd_9[2] .is_wysiwyg = "true";
defparam \rd_9[2] .power_up = "low";

dffeas \rd_10[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[2]~_wirecell_combout ),
	.asdata(\rd_9[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[2]~q ),
	.prn(vcc));
defparam \rd_10[2] .is_wysiwyg = "true";
defparam \rd_10[2] .power_up = "low";

dffeas \rd_11[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[2]~q ),
	.prn(vcc));
defparam \rd_11[2] .is_wysiwyg = "true";
defparam \rd_11[2] .power_up = "low";

dffeas \rd_12[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[2]~q ),
	.prn(vcc));
defparam \rd_12[2] .is_wysiwyg = "true";
defparam \rd_12[2] .power_up = "low";

dffeas \rd_13[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(vcc),
	.asdata(\rd_12[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[2]~q ),
	.prn(vcc));
defparam \rd_13[2] .is_wysiwyg = "true";
defparam \rd_13[2] .power_up = "low";

cyclonev_lcell_comb \rd_14~7 (
	.dataa(!\jam_reg[1]~q ),
	.datab(!\always19~0_combout ),
	.datac(!\rd_14[2]~1_combout ),
	.datad(!\rd_13[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~7 .extended_lut = "off";
defparam \rd_14~7 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \rd_14~7 .shared_arith = "off";

cyclonev_lcell_comb \always19~3_wirecell (
	.dataa(!\always19~3_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always19~3_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always19~3_wirecell .extended_lut = "off";
defparam \always19~3_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \always19~3_wirecell .shared_arith = "off";

dffeas \rd_1[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_7),
	.asdata(dout_reg_sft_31),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[7]~q ),
	.prn(vcc));
defparam \rd_1[7] .is_wysiwyg = "true";
defparam \rd_1[7] .power_up = "low";

dffeas \rd_2[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[7]~q ),
	.prn(vcc));
defparam \rd_2[7] .is_wysiwyg = "true";
defparam \rd_2[7] .power_up = "low";

dffeas \rd_3[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[7]~q ),
	.prn(vcc));
defparam \rd_3[7] .is_wysiwyg = "true";
defparam \rd_3[7] .power_up = "low";

dffeas \rd_4[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[7]~q ),
	.prn(vcc));
defparam \rd_4[7] .is_wysiwyg = "true";
defparam \rd_4[7] .power_up = "low";

dffeas \rd_5[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[7]~q ),
	.prn(vcc));
defparam \rd_5[7] .is_wysiwyg = "true";
defparam \rd_5[7] .power_up = "low";

dffeas \rd_6[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[7]~q ),
	.prn(vcc));
defparam \rd_6[7] .is_wysiwyg = "true";
defparam \rd_6[7] .power_up = "low";

dffeas \rd_7[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[31]~_wirecell_combout ),
	.asdata(\rd_6[7]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[7]~q ),
	.prn(vcc));
defparam \rd_7[7] .is_wysiwyg = "true";
defparam \rd_7[7] .power_up = "low";

dffeas \rd_8[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[23]~_wirecell_combout ),
	.asdata(\rd_7[7]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[7]~q ),
	.prn(vcc));
defparam \rd_8[7] .is_wysiwyg = "true";
defparam \rd_8[7] .power_up = "low";

dffeas \rd_9[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[15]~_wirecell_combout ),
	.asdata(\rd_8[7]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[7]~q ),
	.prn(vcc));
defparam \rd_9[7] .is_wysiwyg = "true";
defparam \rd_9[7] .power_up = "low";

dffeas \rd_10[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[7]~_wirecell_combout ),
	.asdata(\rd_9[7]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[7]~q ),
	.prn(vcc));
defparam \rd_10[7] .is_wysiwyg = "true";
defparam \rd_10[7] .power_up = "low";

dffeas \rd_11[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[7]~q ),
	.prn(vcc));
defparam \rd_11[7] .is_wysiwyg = "true";
defparam \rd_11[7] .power_up = "low";

dffeas \rd_12[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[7]~q ),
	.prn(vcc));
defparam \rd_12[7] .is_wysiwyg = "true";
defparam \rd_12[7] .power_up = "low";

dffeas \rd_13[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always19~3_wirecell_combout ),
	.asdata(\rd_12[7]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[7]~q ),
	.prn(vcc));
defparam \rd_13[7] .is_wysiwyg = "true";
defparam \rd_13[7] .power_up = "low";

cyclonev_lcell_comb \rd_14~8 (
	.dataa(!\jam_reg[2]~q ),
	.datab(!\jam_reg[1]~q ),
	.datac(!\always19~0_combout ),
	.datad(!\rd_14[2]~1_combout ),
	.datae(!\rd_13[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~8 .extended_lut = "off";
defparam \rd_14~8 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \rd_14~8 .shared_arith = "off";

dffeas \rd_1[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(q_b_3),
	.asdata(dout_reg_sft_27),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(!\tx_rden~q ),
	.sload(tx_data_int_7),
	.ena(txclk_ena),
	.q(\rd_1[3]~q ),
	.prn(vcc));
defparam \rd_1[3] .is_wysiwyg = "true";
defparam \rd_1[3] .power_up = "low";

dffeas \rd_2[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_1[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_2[3]~q ),
	.prn(vcc));
defparam \rd_2[3] .is_wysiwyg = "true";
defparam \rd_2[3] .power_up = "low";

dffeas \rd_3[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_2[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_3[3]~q ),
	.prn(vcc));
defparam \rd_3[3] .is_wysiwyg = "true";
defparam \rd_3[3] .power_up = "low";

dffeas \rd_4[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_3[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_4[3]~q ),
	.prn(vcc));
defparam \rd_4[3] .is_wysiwyg = "true";
defparam \rd_4[3] .power_up = "low";

dffeas \rd_5[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_4[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_5[3]~q ),
	.prn(vcc));
defparam \rd_5[3] .is_wysiwyg = "true";
defparam \rd_5[3] .power_up = "low";

dffeas \rd_6[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_5[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_6[3]~q ),
	.prn(vcc));
defparam \rd_6[3] .is_wysiwyg = "true";
defparam \rd_6[3] .power_up = "low";

dffeas \rd_7[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[27]~_wirecell_combout ),
	.asdata(\rd_6[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_7[3]~q ),
	.prn(vcc));
defparam \rd_7[3] .is_wysiwyg = "true";
defparam \rd_7[3] .power_up = "low";

dffeas \rd_8[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[19]~_wirecell_combout ),
	.asdata(\rd_7[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_8[3]~q ),
	.prn(vcc));
defparam \rd_8[3] .is_wysiwyg = "true";
defparam \rd_8[3] .power_up = "low";

dffeas \rd_9[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[11]~_wirecell_combout ),
	.asdata(\rd_8[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_9[3]~q ),
	.prn(vcc));
defparam \rd_9[3] .is_wysiwyg = "true";
defparam \rd_9[3] .power_up = "low";

dffeas \rd_10[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_CRC|U_GALS|reg_out[3]~_wirecell_combout ),
	.asdata(\rd_9[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always17~1_combout ),
	.ena(txclk_ena),
	.q(\rd_10[3]~q ),
	.prn(vcc));
defparam \rd_10[3] .is_wysiwyg = "true";
defparam \rd_10[3] .power_up = "low";

dffeas \rd_11[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_10[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_11[3]~q ),
	.prn(vcc));
defparam \rd_11[3] .is_wysiwyg = "true";
defparam \rd_11[3] .power_up = "low";

dffeas \rd_12[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\rd_11[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\rd_12[3]~q ),
	.prn(vcc));
defparam \rd_12[3] .is_wysiwyg = "true";
defparam \rd_12[3] .power_up = "low";

dffeas \rd_13[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(GND_port),
	.asdata(\rd_12[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\always19~1_combout ),
	.sload(\rd_13[6]~0_combout ),
	.ena(txclk_ena),
	.q(\rd_13[3]~q ),
	.prn(vcc));
defparam \rd_13[3] .is_wysiwyg = "true";
defparam \rd_13[3] .power_up = "low";

cyclonev_lcell_comb \rd_14~9 (
	.dataa(!\rd_14[2]~1_combout ),
	.datab(!\rd_13[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rd_14~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rd_14~9 .extended_lut = "off";
defparam \rd_14~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \rd_14~9 .shared_arith = "off";

cyclonev_lcell_comb \always14~0 (
	.dataa(!\tx_rden~q ),
	.datab(!empty_flag),
	.datac(!tx_stat_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~0 .extended_lut = "off";
defparam \always14~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always14~0 .shared_arith = "off";

dffeas \tx_err_s[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\always14~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[0]~q ),
	.prn(vcc));
defparam \tx_err_s[0] .is_wysiwyg = "true";
defparam \tx_err_s[0] .power_up = "low";

dffeas \tx_err_s[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[1]~q ),
	.prn(vcc));
defparam \tx_err_s[1] .is_wysiwyg = "true";
defparam \tx_err_s[1] .power_up = "low";

cyclonev_lcell_comb \tx_err_s~0 (
	.dataa(!\frm_rd[2]~q ),
	.datab(!\tx_err_s[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_err_s~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_err_s~0 .extended_lut = "off";
defparam \tx_err_s~0 .lut_mask = 64'h7777777777777777;
defparam \tx_err_s~0 .shared_arith = "off";

dffeas \tx_err_s[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[2]~q ),
	.prn(vcc));
defparam \tx_err_s[2] .is_wysiwyg = "true";
defparam \tx_err_s[2] .power_up = "low";

dffeas \tx_err_s[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[3]~q ),
	.prn(vcc));
defparam \tx_err_s[3] .is_wysiwyg = "true";
defparam \tx_err_s[3] .power_up = "low";

dffeas \tx_err_s[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_err_s[4]~q ),
	.prn(vcc));
defparam \tx_err_s[4] .is_wysiwyg = "true";
defparam \tx_err_s[4] .power_up = "low";

dffeas \tx_err_s[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[5]~q ),
	.prn(vcc));
defparam \tx_err_s[5] .is_wysiwyg = "true";
defparam \tx_err_s[5] .power_up = "low";

dffeas \tx_err_s[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[6]~q ),
	.prn(vcc));
defparam \tx_err_s[6] .is_wysiwyg = "true";
defparam \tx_err_s[6] .power_up = "low";

dffeas \tx_err_s[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[7]~q ),
	.prn(vcc));
defparam \tx_err_s[7] .is_wysiwyg = "true";
defparam \tx_err_s[7] .power_up = "low";

dffeas \tx_err_s[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[7]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[8]~q ),
	.prn(vcc));
defparam \tx_err_s[8] .is_wysiwyg = "true";
defparam \tx_err_s[8] .power_up = "low";

dffeas \tx_err_s[9] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[8]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[9]~q ),
	.prn(vcc));
defparam \tx_err_s[9] .is_wysiwyg = "true";
defparam \tx_err_s[9] .power_up = "low";

dffeas \tx_err_s[10] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[9]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[10]~q ),
	.prn(vcc));
defparam \tx_err_s[10] .is_wysiwyg = "true";
defparam \tx_err_s[10] .power_up = "low";

dffeas \tx_err_s[11] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[10]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[11]~q ),
	.prn(vcc));
defparam \tx_err_s[11] .is_wysiwyg = "true";
defparam \tx_err_s[11] .power_up = "low";

dffeas \tx_err_s[12] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[11]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[12]~q ),
	.prn(vcc));
defparam \tx_err_s[12] .is_wysiwyg = "true";
defparam \tx_err_s[12] .power_up = "low";

dffeas \tx_err_s[13] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[12]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[13]~q ),
	.prn(vcc));
defparam \tx_err_s[13] .is_wysiwyg = "true";
defparam \tx_err_s[13] .power_up = "low";

dffeas \tx_err_s[14] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[13]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[14]~q ),
	.prn(vcc));
defparam \tx_err_s[14] .is_wysiwyg = "true";
defparam \tx_err_s[14] .power_up = "low";

dffeas \tx_err_s[15] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[14]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[15]~q ),
	.prn(vcc));
defparam \tx_err_s[15] .is_wysiwyg = "true";
defparam \tx_err_s[15] .power_up = "low";

dffeas \tx_err_s[16] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[15]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[16]~q ),
	.prn(vcc));
defparam \tx_err_s[16] .is_wysiwyg = "true";
defparam \tx_err_s[16] .power_up = "low";

dffeas \tx_err_s[17] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[16]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[17]~q ),
	.prn(vcc));
defparam \tx_err_s[17] .is_wysiwyg = "true";
defparam \tx_err_s[17] .power_up = "low";

dffeas \tx_err_s[18] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[17]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[18]~q ),
	.prn(vcc));
defparam \tx_err_s[18] .is_wysiwyg = "true";
defparam \tx_err_s[18] .power_up = "low";

dffeas \tx_err_s[19] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_err_s[18]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_err_s[19]~q ),
	.prn(vcc));
defparam \tx_err_s[19] .is_wysiwyg = "true";
defparam \tx_err_s[19] .power_up = "low";

cyclonev_lcell_comb \tx_err~0 (
	.dataa(!\tx_err_s[19]~q ),
	.datab(!\tx_err_s[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_err~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_err~0 .extended_lut = "off";
defparam \tx_err~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \tx_err~0 .shared_arith = "off";

cyclonev_lcell_comb \gm_rx_crs_reg3~0 (
	.dataa(!\gap_wait~q ),
	.datab(!dreg_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gm_rx_crs_reg3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gm_rx_crs_reg3~0 .extended_lut = "off";
defparam \gm_rx_crs_reg3~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \gm_rx_crs_reg3~0 .shared_arith = "off";

dffeas gm_rx_crs_reg3(
	.clk(mac_tx_clock_connection_clk),
	.d(\gm_rx_crs_reg3~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gm_rx_crs_reg3~q ),
	.prn(vcc));
defparam gm_rx_crs_reg3.is_wysiwyg = "true";
defparam gm_rx_crs_reg3.power_up = "low";

cyclonev_lcell_comb \gm_rx_crs_reg4~0 (
	.dataa(!\gap_wait~q ),
	.datab(!\gm_rx_crs_reg3~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gm_rx_crs_reg4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gm_rx_crs_reg4~0 .extended_lut = "off";
defparam \gm_rx_crs_reg4~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \gm_rx_crs_reg4~0 .shared_arith = "off";

dffeas gm_rx_crs_reg4(
	.clk(mac_tx_clock_connection_clk),
	.d(\gm_rx_crs_reg4~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\gm_rx_crs_reg4~q ),
	.prn(vcc));
defparam gm_rx_crs_reg4.is_wysiwyg = "true";
defparam gm_rx_crs_reg4.power_up = "low";

cyclonev_lcell_comb \frm_wait~0 (
	.dataa(!dreg_1),
	.datab(!\gm_rx_col_reg2~q ),
	.datac(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datad(!col_int1),
	.datae(!\gm_rx_crs_reg4~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_wait~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_wait~0 .extended_lut = "off";
defparam \frm_wait~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \frm_wait~0 .shared_arith = "off";

dffeas tx_sav_int_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(tx_sav_int),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_sav_int_reg~q ),
	.prn(vcc));
defparam tx_sav_int_reg.is_wysiwyg = "true";
defparam tx_sav_int_reg.power_up = "low";

cyclonev_lcell_comb \frm_wait~1 (
	.dataa(!\frm_wait~q ),
	.datab(!\gap_wait~q ),
	.datac(!\tx_sav_int_reg~q ),
	.datad(!empty_flag),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_wait~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_wait~1 .extended_lut = "off";
defparam \frm_wait~1 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \frm_wait~1 .shared_arith = "off";

cyclonev_lcell_comb \frm_wait~2 (
	.dataa(!\frm_rd[2]~q ),
	.datab(!\U_SYNC_MAGIC_ENA|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_SLEEP_ENA|std_sync_no_cut|dreg[1]~q ),
	.datad(!\frm_rd[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_wait~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_wait~2 .extended_lut = "off";
defparam \frm_wait~2 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \frm_wait~2 .shared_arith = "off";

cyclonev_lcell_comb \frm_wait~3 (
	.dataa(!\U_SYNC_2|std_sync_no_cut|dreg[1]~q ),
	.datab(!mac_ena),
	.datac(!\frm_wait~0_combout ),
	.datad(!\frm_wait~1_combout ),
	.datae(!\frm_wait~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\frm_wait~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \frm_wait~3 .extended_lut = "off";
defparam \frm_wait~3 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \frm_wait~3 .shared_arith = "off";

dffeas frm_wait(
	.clk(mac_tx_clock_connection_clk),
	.d(\frm_wait~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\frm_wait~q ),
	.prn(vcc));
defparam frm_wait.is_wysiwyg = "true";
defparam frm_wait.power_up = "low";

dffeas \tx_en_s[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(tx_en_s_1),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_en_s[2]~q ),
	.prn(vcc));
defparam \tx_en_s[2] .is_wysiwyg = "true";
defparam \tx_en_s[2] .power_up = "low";

dffeas \tx_en_s[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\tx_en_s[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(txclk_ena),
	.q(\tx_en_s[3]~q ),
	.prn(vcc));
defparam \tx_en_s[3] .is_wysiwyg = "true";
defparam \tx_en_s[3] .power_up = "low";

cyclonev_lcell_comb \col_int~0 (
	.dataa(!dreg_1),
	.datab(!tx_en_s_1),
	.datac(!\gm_rx_col_reg2~q ),
	.datad(!\U_SYNC_4|std_sync_no_cut|dreg[1]~q ),
	.datae(!col_int1),
	.dataf(!\tx_en_s[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\col_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_int~0 .extended_lut = "off";
defparam \col_int~0 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \col_int~0 .shared_arith = "off";

cyclonev_lcell_comb \always9~5 (
	.dataa(!txclk_ena),
	.datab(!\always9~0_combout ),
	.datac(!\eop_0~1_combout ),
	.datad(!always9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~5 .extended_lut = "off";
defparam \always9~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \always9~5 .shared_arith = "off";

cyclonev_lcell_comb \always6~3 (
	.dataa(!txclk_ena),
	.datab(!\frm_rd[0]~q ),
	.datac(!\eop_0~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~3 .extended_lut = "off";
defparam \always6~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always6~3 .shared_arith = "off";

dffeas tx_stat_rden_i(
	.clk(mac_tx_clock_connection_clk),
	.d(\always6~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tx_stat_rden_i~q ),
	.prn(vcc));
defparam tx_stat_rden_i.is_wysiwyg = "true";
defparam tx_stat_rden_i.power_up = "low";

cyclonev_lcell_comb \tx_stat_rden~0 (
	.dataa(!\always3~0_combout ),
	.datab(!\tx_stat_rden_i~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_stat_rden~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_stat_rden~0 .extended_lut = "off";
defparam \tx_stat_rden~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \tx_stat_rden~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_128 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	ethernet_mode,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	ethernet_mode;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_128 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(ethernet_mode),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_128 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_129 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_129 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_129 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_130 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_130 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_130 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_131 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	m_rx_crs,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	m_rx_crs;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_131 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(m_rx_crs),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_131 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_132 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	gm_rx_col_reg,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	gm_rx_col_reg;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_132 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(gm_rx_col_reg),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_132 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_133 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_133 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_133 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_134 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	sleep_ena,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	sleep_ena;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_134 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(sleep_ena),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_134 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_9 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_139 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_138 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_137 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_136 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_135 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_135 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_135 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_135 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_136 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_136 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_136 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_137 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_137 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_137 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_138 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_138 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_138 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_139 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_139 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_139 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_crc328generator (
	txclk_ena,
	altera_tse_reset_synchronizer_chain_out,
	sop_4,
	eof_dly_5,
	rd_5_4,
	rd_5_0,
	rd_5_5,
	rd_5_1,
	rd_5_6,
	rd_5_2,
	rd_5_7,
	rd_5_3,
	eop_4,
	reg_out_0,
	reg_out_10,
	reg_out_11,
	reg_out_12,
	reg_out_13,
	reg_out_14,
	reg_out_15,
	reg_out_16,
	reg_out_17,
	reg_out_18,
	reg_out_19,
	reg_out_1,
	reg_out_20,
	reg_out_21,
	reg_out_22,
	reg_out_23,
	reg_out_24,
	reg_out_25,
	reg_out_26,
	reg_out_27,
	reg_out_28,
	reg_out_29,
	reg_out_2,
	reg_out_30,
	reg_out_31,
	reg_out_3,
	reg_out_4,
	reg_out_5,
	reg_out_6,
	reg_out_7,
	reg_out_8,
	reg_out_9,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	txclk_ena;
input 	altera_tse_reset_synchronizer_chain_out;
input 	sop_4;
output 	eof_dly_5;
input 	rd_5_4;
input 	rd_5_0;
input 	rd_5_5;
input 	rd_5_1;
input 	rd_5_6;
input 	rd_5_2;
input 	rd_5_7;
input 	rd_5_3;
input 	eop_4;
output 	reg_out_0;
output 	reg_out_10;
output 	reg_out_11;
output 	reg_out_12;
output 	reg_out_13;
output 	reg_out_14;
output 	reg_out_15;
output 	reg_out_16;
output 	reg_out_17;
output 	reg_out_18;
output 	reg_out_19;
output 	reg_out_1;
output 	reg_out_20;
output 	reg_out_21;
output 	reg_out_22;
output 	reg_out_23;
output 	reg_out_24;
output 	reg_out_25;
output 	reg_out_26;
output 	reg_out_27;
output 	reg_out_28;
output 	reg_out_29;
output 	reg_out_2;
output 	reg_out_30;
output 	reg_out_31;
output 	reg_out_3;
output 	reg_out_4;
output 	reg_out_5;
output 	reg_out_6;
output 	reg_out_7;
output 	reg_out_8;
output 	reg_out_9;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_tse_crc32ctl8 U_CTL(
	.clk_ena(txclk_ena),
	.rst(altera_tse_reset_synchronizer_chain_out),
	.eof_dly_5(eof_dly_5),
	.eof(eop_4),
	.clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_crc32galois8_1 U_GALS(
	.clk_ena(txclk_ena),
	.rst(altera_tse_reset_synchronizer_chain_out),
	.sop_4(sop_4),
	.rd_5_4(rd_5_4),
	.rd_5_0(rd_5_0),
	.rd_5_5(rd_5_5),
	.rd_5_1(rd_5_1),
	.rd_5_6(rd_5_6),
	.rd_5_2(rd_5_2),
	.rd_5_7(rd_5_7),
	.rd_5_3(rd_5_3),
	.reg_out_0(reg_out_0),
	.reg_out_10(reg_out_10),
	.reg_out_11(reg_out_11),
	.reg_out_12(reg_out_12),
	.reg_out_13(reg_out_13),
	.reg_out_14(reg_out_14),
	.reg_out_15(reg_out_15),
	.reg_out_16(reg_out_16),
	.reg_out_17(reg_out_17),
	.reg_out_18(reg_out_18),
	.reg_out_19(reg_out_19),
	.reg_out_1(reg_out_1),
	.reg_out_20(reg_out_20),
	.reg_out_21(reg_out_21),
	.reg_out_22(reg_out_22),
	.reg_out_23(reg_out_23),
	.reg_out_24(reg_out_24),
	.reg_out_25(reg_out_25),
	.reg_out_26(reg_out_26),
	.reg_out_27(reg_out_27),
	.reg_out_28(reg_out_28),
	.reg_out_29(reg_out_29),
	.reg_out_2(reg_out_2),
	.reg_out_30(reg_out_30),
	.reg_out_31(reg_out_31),
	.reg_out_3(reg_out_3),
	.reg_out_4(reg_out_4),
	.reg_out_5(reg_out_5),
	.reg_out_6(reg_out_6),
	.reg_out_7(reg_out_7),
	.reg_out_8(reg_out_8),
	.reg_out_9(reg_out_9),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_tse_crc32ctl8 (
	clk_ena,
	rst,
	eof_dly_5,
	eof,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clk_ena;
input 	rst;
output 	eof_dly_5;
input 	eof;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \eof_dly[0]~q ;
wire \eof_dly[1]~q ;
wire \eof_dly[2]~q ;
wire \eof_dly[3]~q ;
wire \eof_dly[4]~q ;


dffeas \eof_dly[5] (
	.clk(clk),
	.d(\eof_dly[4]~q ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(eof_dly_5),
	.prn(vcc));
defparam \eof_dly[5] .is_wysiwyg = "true";
defparam \eof_dly[5] .power_up = "low";

dffeas \eof_dly[0] (
	.clk(clk),
	.d(eof),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\eof_dly[0]~q ),
	.prn(vcc));
defparam \eof_dly[0] .is_wysiwyg = "true";
defparam \eof_dly[0] .power_up = "low";

dffeas \eof_dly[1] (
	.clk(clk),
	.d(\eof_dly[0]~q ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\eof_dly[1]~q ),
	.prn(vcc));
defparam \eof_dly[1] .is_wysiwyg = "true";
defparam \eof_dly[1] .power_up = "low";

dffeas \eof_dly[2] (
	.clk(clk),
	.d(\eof_dly[1]~q ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\eof_dly[2]~q ),
	.prn(vcc));
defparam \eof_dly[2] .is_wysiwyg = "true";
defparam \eof_dly[2] .power_up = "low";

dffeas \eof_dly[3] (
	.clk(clk),
	.d(\eof_dly[2]~q ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\eof_dly[3]~q ),
	.prn(vcc));
defparam \eof_dly[3] .is_wysiwyg = "true";
defparam \eof_dly[3] .power_up = "low";

dffeas \eof_dly[4] (
	.clk(clk),
	.d(\eof_dly[3]~q ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\eof_dly[4]~q ),
	.prn(vcc));
defparam \eof_dly[4] .is_wysiwyg = "true";
defparam \eof_dly[4] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_crc32galois8_1 (
	clk_ena,
	rst,
	sop_4,
	rd_5_4,
	rd_5_0,
	rd_5_5,
	rd_5_1,
	rd_5_6,
	rd_5_2,
	rd_5_7,
	rd_5_3,
	reg_out_0,
	reg_out_10,
	reg_out_11,
	reg_out_12,
	reg_out_13,
	reg_out_14,
	reg_out_15,
	reg_out_16,
	reg_out_17,
	reg_out_18,
	reg_out_19,
	reg_out_1,
	reg_out_20,
	reg_out_21,
	reg_out_22,
	reg_out_23,
	reg_out_24,
	reg_out_25,
	reg_out_26,
	reg_out_27,
	reg_out_28,
	reg_out_29,
	reg_out_2,
	reg_out_30,
	reg_out_31,
	reg_out_3,
	reg_out_4,
	reg_out_5,
	reg_out_6,
	reg_out_7,
	reg_out_8,
	reg_out_9,
	clk)/* synthesis synthesis_greybox=1 */;
input 	clk_ena;
input 	rst;
input 	sop_4;
input 	rd_5_4;
input 	rd_5_0;
input 	rd_5_5;
input 	rd_5_1;
input 	rd_5_6;
input 	rd_5_2;
input 	rd_5_7;
input 	rd_5_3;
output 	reg_out_0;
output 	reg_out_10;
output 	reg_out_11;
output 	reg_out_12;
output 	reg_out_13;
output 	reg_out_14;
output 	reg_out_15;
output 	reg_out_16;
output 	reg_out_17;
output 	reg_out_18;
output 	reg_out_19;
output 	reg_out_1;
output 	reg_out_20;
output 	reg_out_21;
output 	reg_out_22;
output 	reg_out_23;
output 	reg_out_24;
output 	reg_out_25;
output 	reg_out_26;
output 	reg_out_27;
output 	reg_out_28;
output 	reg_out_29;
output 	reg_out_2;
output 	reg_out_30;
output 	reg_out_31;
output 	reg_out_3;
output 	reg_out_4;
output 	reg_out_5;
output 	reg_out_6;
output 	reg_out_7;
output 	reg_out_8;
output 	reg_out_9;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \o[31]~combout ;
wire \reg_out[31]~q ;
wire \o[23]~combout ;
wire \reg_out[23]~q ;
wire \o[15]~combout ;
wire \reg_out[15]~q ;
wire \o[7]~combout ;
wire \reg_out[7]~q ;
wire \o[27]~combout ;
wire \reg_out[27]~q ;
wire \o[19]~1_combout ;
wire \o[19]~combout ;
wire \reg_out[19]~q ;
wire \o[11]~combout ;
wire \reg_out[11]~q ;
wire \o[3]~combout ;
wire \reg_out[3]~q ;
wire \o1[17]~0_combout ;
wire \o[25]~combout ;
wire \reg_out[25]~q ;
wire \o[17]~combout ;
wire \reg_out[17]~q ;
wire \o[9]~combout ;
wire \reg_out[9]~q ;
wire \o[1]~combout ;
wire \reg_out[1]~q ;
wire \o[29]~combout ;
wire \reg_out[29]~q ;
wire \o[21]~combout ;
wire \reg_out[21]~q ;
wire \o[13]~combout ;
wire \reg_out[13]~q ;
wire \o[5]~combout ;
wire \reg_out[5]~q ;
wire \o[30]~combout ;
wire \reg_out[30]~q ;
wire \o[22]~combout ;
wire \reg_out[22]~q ;
wire \o[14]~combout ;
wire \reg_out[14]~q ;
wire \o[6]~combout ;
wire \reg_out[6]~q ;
wire \o1[0]~combout ;
wire \o[28]~combout ;
wire \reg_out[28]~q ;
wire \o[20]~combout ;
wire \reg_out[20]~q ;
wire \o[12]~combout ;
wire \reg_out[12]~q ;
wire \o[4]~combout ;
wire \reg_out[4]~q ;
wire \o[26]~combout ;
wire \reg_out[26]~q ;
wire \o[18]~0_combout ;
wire \o[18]~combout ;
wire \reg_out[18]~q ;
wire \o[10]~combout ;
wire \reg_out[10]~q ;
wire \o[2]~combout ;
wire \reg_out[2]~q ;
wire \o[24]~combout ;
wire \reg_out[24]~q ;
wire \o[16]~combout ;
wire \reg_out[16]~q ;
wire \o[8]~combout ;
wire \reg_out[8]~q ;
wire \o[0]~combout ;
wire \reg_out[0]~q ;


cyclonev_lcell_comb \reg_out[0]~_wirecell (
	.dataa(!\reg_out[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[0]~_wirecell .extended_lut = "off";
defparam \reg_out[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[0]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[10]~_wirecell (
	.dataa(!\reg_out[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[10]~_wirecell .extended_lut = "off";
defparam \reg_out[10]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[10]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[11]~_wirecell (
	.dataa(!\reg_out[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[11]~_wirecell .extended_lut = "off";
defparam \reg_out[11]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[11]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[12]~_wirecell (
	.dataa(!\reg_out[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[12]~_wirecell .extended_lut = "off";
defparam \reg_out[12]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[12]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[13]~_wirecell (
	.dataa(!\reg_out[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[13]~_wirecell .extended_lut = "off";
defparam \reg_out[13]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[13]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[14]~_wirecell (
	.dataa(!\reg_out[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[14]~_wirecell .extended_lut = "off";
defparam \reg_out[14]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[14]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[15]~_wirecell (
	.dataa(!\reg_out[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[15]~_wirecell .extended_lut = "off";
defparam \reg_out[15]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[15]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[16]~_wirecell (
	.dataa(!\reg_out[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[16]~_wirecell .extended_lut = "off";
defparam \reg_out[16]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[16]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[17]~_wirecell (
	.dataa(!\reg_out[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[17]~_wirecell .extended_lut = "off";
defparam \reg_out[17]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[17]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[18]~_wirecell (
	.dataa(!\reg_out[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[18]~_wirecell .extended_lut = "off";
defparam \reg_out[18]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[18]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[19]~_wirecell (
	.dataa(!\reg_out[19]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[19]~_wirecell .extended_lut = "off";
defparam \reg_out[19]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[19]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[1]~_wirecell (
	.dataa(!\reg_out[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[1]~_wirecell .extended_lut = "off";
defparam \reg_out[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[20]~_wirecell (
	.dataa(!\reg_out[20]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[20]~_wirecell .extended_lut = "off";
defparam \reg_out[20]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[20]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[21]~_wirecell (
	.dataa(!\reg_out[21]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[21]~_wirecell .extended_lut = "off";
defparam \reg_out[21]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[21]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[22]~_wirecell (
	.dataa(!\reg_out[22]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[22]~_wirecell .extended_lut = "off";
defparam \reg_out[22]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[22]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[23]~_wirecell (
	.dataa(!\reg_out[23]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[23]~_wirecell .extended_lut = "off";
defparam \reg_out[23]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[23]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[24]~_wirecell (
	.dataa(!\reg_out[24]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[24]~_wirecell .extended_lut = "off";
defparam \reg_out[24]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[24]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[25]~_wirecell (
	.dataa(!\reg_out[25]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[25]~_wirecell .extended_lut = "off";
defparam \reg_out[25]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[25]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[26]~_wirecell (
	.dataa(!\reg_out[26]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[26]~_wirecell .extended_lut = "off";
defparam \reg_out[26]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[26]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[27]~_wirecell (
	.dataa(!\reg_out[27]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[27]~_wirecell .extended_lut = "off";
defparam \reg_out[27]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[27]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[28]~_wirecell (
	.dataa(!\reg_out[28]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[28]~_wirecell .extended_lut = "off";
defparam \reg_out[28]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[28]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[29]~_wirecell (
	.dataa(!\reg_out[29]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[29]~_wirecell .extended_lut = "off";
defparam \reg_out[29]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[29]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[2]~_wirecell (
	.dataa(!\reg_out[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[2]~_wirecell .extended_lut = "off";
defparam \reg_out[2]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[2]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[30]~_wirecell (
	.dataa(!\reg_out[30]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[30]~_wirecell .extended_lut = "off";
defparam \reg_out[30]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[30]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[31]~_wirecell (
	.dataa(!\reg_out[31]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[31]~_wirecell .extended_lut = "off";
defparam \reg_out[31]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[31]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[3]~_wirecell (
	.dataa(!\reg_out[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[3]~_wirecell .extended_lut = "off";
defparam \reg_out[3]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[3]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[4]~_wirecell (
	.dataa(!\reg_out[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[4]~_wirecell .extended_lut = "off";
defparam \reg_out[4]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[4]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[5]~_wirecell (
	.dataa(!\reg_out[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[5]~_wirecell .extended_lut = "off";
defparam \reg_out[5]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[5]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[6]~_wirecell (
	.dataa(!\reg_out[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[6]~_wirecell .extended_lut = "off";
defparam \reg_out[6]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[6]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[7]~_wirecell (
	.dataa(!\reg_out[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[7]~_wirecell .extended_lut = "off";
defparam \reg_out[7]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[7]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[8]~_wirecell (
	.dataa(!\reg_out[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[8]~_wirecell .extended_lut = "off";
defparam \reg_out[8]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[8]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \reg_out[9]~_wirecell (
	.dataa(!\reg_out[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(reg_out_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \reg_out[9]~_wirecell .extended_lut = "off";
defparam \reg_out[9]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \reg_out[9]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \o[31] (
	.dataa(!\reg_out[1]~q ),
	.datab(!\reg_out[7]~q ),
	.datac(!rd_5_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[31] .extended_lut = "off";
defparam \o[31] .lut_mask = 64'h9696969696969696;
defparam \o[31] .shared_arith = "off";

dffeas \reg_out[31] (
	.clk(clk),
	.d(\o[31]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[31]~q ),
	.prn(vcc));
defparam \reg_out[31] .is_wysiwyg = "true";
defparam \reg_out[31] .power_up = "low";

cyclonev_lcell_comb \o[23] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[7]~q ),
	.datad(!\reg_out[3]~q ),
	.datae(!\reg_out[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[23] .extended_lut = "off";
defparam \o[23] .lut_mask = 64'h9669699696696996;
defparam \o[23] .shared_arith = "off";

dffeas \reg_out[23] (
	.clk(clk),
	.d(\o[23]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[23]~q ),
	.prn(vcc));
defparam \reg_out[23] .is_wysiwyg = "true";
defparam \reg_out[23] .power_up = "low";

cyclonev_lcell_comb \o[15] (
	.dataa(!\reg_out[2]~q ),
	.datab(!\reg_out[7]~q ),
	.datac(!\reg_out[3]~q ),
	.datad(!\reg_out[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[15] .extended_lut = "off";
defparam \o[15] .lut_mask = 64'h6996699669966996;
defparam \o[15] .shared_arith = "off";

dffeas \reg_out[15] (
	.clk(clk),
	.d(\o[15]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[15]~q ),
	.prn(vcc));
defparam \reg_out[15] .is_wysiwyg = "true";
defparam \reg_out[15] .power_up = "low";

cyclonev_lcell_comb \o[7] (
	.dataa(!\reg_out[0]~q ),
	.datab(!\reg_out[5]~q ),
	.datac(!\reg_out[6]~q ),
	.datad(!\reg_out[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[7] .extended_lut = "off";
defparam \o[7] .lut_mask = 64'h6996699669966996;
defparam \o[7] .shared_arith = "off";

dffeas \reg_out[7] (
	.clk(clk),
	.d(\o[7]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[7]~q ),
	.prn(vcc));
defparam \reg_out[7] .is_wysiwyg = "true";
defparam \reg_out[7] .power_up = "low";

cyclonev_lcell_comb \o[27] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[5]~q ),
	.datac(!\reg_out[1]~q ),
	.datad(!\reg_out[7]~q ),
	.datae(!\reg_out[3]~q ),
	.dataf(!rd_5_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[27] .extended_lut = "off";
defparam \o[27] .lut_mask = 64'h6996966996696996;
defparam \o[27] .shared_arith = "off";

dffeas \reg_out[27] (
	.clk(clk),
	.d(\o[27]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[27]~q ),
	.prn(vcc));
defparam \reg_out[27] .is_wysiwyg = "true";
defparam \reg_out[27] .power_up = "low";

cyclonev_lcell_comb \o[19]~1 (
	.dataa(!\reg_out[6]~q ),
	.datab(!\reg_out[7]~q ),
	.datac(!\reg_out[3]~q ),
	.datad(!\reg_out[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[19]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[19]~1 .extended_lut = "off";
defparam \o[19]~1 .lut_mask = 64'h6996699669966996;
defparam \o[19]~1 .shared_arith = "off";

cyclonev_lcell_comb \o[19] (
	.dataa(!\reg_out[5]~q ),
	.datab(!\reg_out[1]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\o[19]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[19] .extended_lut = "off";
defparam \o[19] .lut_mask = 64'h6996699669966996;
defparam \o[19] .shared_arith = "off";

dffeas \reg_out[19] (
	.clk(clk),
	.d(\o[19]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[19]~q ),
	.prn(vcc));
defparam \reg_out[19] .is_wysiwyg = "true";
defparam \reg_out[19] .power_up = "low";

cyclonev_lcell_comb \o[11] (
	.dataa(!\reg_out[3]~q ),
	.datab(!\reg_out[19]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[11] .extended_lut = "off";
defparam \o[11] .lut_mask = 64'h6666666666666666;
defparam \o[11] .shared_arith = "off";

dffeas \reg_out[11] (
	.clk(clk),
	.d(\o[11]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[11]~q ),
	.prn(vcc));
defparam \reg_out[11] .is_wysiwyg = "true";
defparam \reg_out[11] .power_up = "low";

cyclonev_lcell_comb \o[3] (
	.dataa(!\reg_out[5]~q ),
	.datab(!\reg_out[1]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[3] .extended_lut = "off";
defparam \o[3] .lut_mask = 64'h6996699669966996;
defparam \o[3] .shared_arith = "off";

dffeas \reg_out[3] (
	.clk(clk),
	.d(\o[3]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[3]~q ),
	.prn(vcc));
defparam \reg_out[3] .is_wysiwyg = "true";
defparam \reg_out[3] .power_up = "low";

cyclonev_lcell_comb \o1[17]~0 (
	.dataa(!\reg_out[0]~q ),
	.datab(!\reg_out[5]~q ),
	.datac(!\reg_out[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o1[17]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o1[17]~0 .extended_lut = "off";
defparam \o1[17]~0 .lut_mask = 64'h9696969696969696;
defparam \o1[17]~0 .shared_arith = "off";

cyclonev_lcell_comb \o[25] (
	.dataa(!\reg_out[5]~q ),
	.datab(!\reg_out[1]~q ),
	.datac(!\o1[0]~combout ),
	.datad(!rd_5_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[25] .extended_lut = "off";
defparam \o[25] .lut_mask = 64'h6996699669966996;
defparam \o[25] .shared_arith = "off";

dffeas \reg_out[25] (
	.clk(clk),
	.d(\o[25]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[25]~q ),
	.prn(vcc));
defparam \reg_out[25] .is_wysiwyg = "true";
defparam \reg_out[25] .power_up = "low";

cyclonev_lcell_comb \o[17] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[3]~q ),
	.datac(!\o1[17]~0_combout ),
	.datad(!\reg_out[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[17] .extended_lut = "off";
defparam \o[17] .lut_mask = 64'h6996699669966996;
defparam \o[17] .shared_arith = "off";

dffeas \reg_out[17] (
	.clk(clk),
	.d(\o[17]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[17]~q ),
	.prn(vcc));
defparam \reg_out[17] .is_wysiwyg = "true";
defparam \reg_out[17] .power_up = "low";

cyclonev_lcell_comb \o[9] (
	.dataa(!\reg_out[7]~q ),
	.datab(!\reg_out[17]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[9] .extended_lut = "off";
defparam \o[9] .lut_mask = 64'h6666666666666666;
defparam \o[9] .shared_arith = "off";

dffeas \reg_out[9] (
	.clk(clk),
	.d(\o[9]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[9]~q ),
	.prn(vcc));
defparam \reg_out[9] .is_wysiwyg = "true";
defparam \reg_out[9] .power_up = "low";

cyclonev_lcell_comb \o[1] (
	.dataa(!\reg_out[0]~q ),
	.datab(!\reg_out[3]~q ),
	.datac(!\reg_out[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[1] .extended_lut = "off";
defparam \o[1] .lut_mask = 64'h9696969696969696;
defparam \o[1] .shared_arith = "off";

dffeas \reg_out[1] (
	.clk(clk),
	.d(\o[1]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[1]~q ),
	.prn(vcc));
defparam \reg_out[1] .is_wysiwyg = "true";
defparam \reg_out[1] .power_up = "low";

cyclonev_lcell_comb \o[29] (
	.dataa(!\reg_out[6]~q ),
	.datab(!\reg_out[7]~q ),
	.datac(!\o1[17]~0_combout ),
	.datad(!rd_5_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[29] .extended_lut = "off";
defparam \o[29] .lut_mask = 64'h6996699669966996;
defparam \o[29] .shared_arith = "off";

dffeas \reg_out[29] (
	.clk(clk),
	.d(\o[29]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[29]~q ),
	.prn(vcc));
defparam \reg_out[29] .is_wysiwyg = "true";
defparam \reg_out[29] .power_up = "low";

cyclonev_lcell_comb \o[21] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[5]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[7]~q ),
	.datae(!\reg_out[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[21] .extended_lut = "off";
defparam \o[21] .lut_mask = 64'h9669699696696996;
defparam \o[21] .shared_arith = "off";

dffeas \reg_out[21] (
	.clk(clk),
	.d(\o[21]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[21]~q ),
	.prn(vcc));
defparam \reg_out[21] .is_wysiwyg = "true";
defparam \reg_out[21] .power_up = "low";

cyclonev_lcell_comb \o[13] (
	.dataa(!\reg_out[21]~q ),
	.datab(!\o1[17]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[13] .extended_lut = "off";
defparam \o[13] .lut_mask = 64'h6666666666666666;
defparam \o[13] .shared_arith = "off";

dffeas \reg_out[13] (
	.clk(clk),
	.d(\o[13]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[13]~q ),
	.prn(vcc));
defparam \reg_out[13] .is_wysiwyg = "true";
defparam \reg_out[13] .power_up = "low";

cyclonev_lcell_comb \o[5] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[1]~q ),
	.datac(!\reg_out[7]~q ),
	.datad(!\reg_out[3]~q ),
	.datae(!\reg_out[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[5] .extended_lut = "off";
defparam \o[5] .lut_mask = 64'h9669699696696996;
defparam \o[5] .shared_arith = "off";

dffeas \reg_out[5] (
	.clk(clk),
	.d(\o[5]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[5]~q ),
	.prn(vcc));
defparam \reg_out[5] .is_wysiwyg = "true";
defparam \reg_out[5] .power_up = "low";

cyclonev_lcell_comb \o[30] (
	.dataa(!\reg_out[0]~q ),
	.datab(!\reg_out[1]~q ),
	.datac(!\reg_out[6]~q ),
	.datad(!\reg_out[7]~q ),
	.datae(!rd_5_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[30] .extended_lut = "off";
defparam \o[30] .lut_mask = 64'h9669699696696996;
defparam \o[30] .shared_arith = "off";

dffeas \reg_out[30] (
	.clk(clk),
	.d(\o[30]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[30]~q ),
	.prn(vcc));
defparam \reg_out[30] .is_wysiwyg = "true";
defparam \reg_out[30] .power_up = "low";

cyclonev_lcell_comb \o[22] (
	.dataa(!\reg_out[5]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[3]~q ),
	.datae(!\reg_out[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[22] .extended_lut = "off";
defparam \o[22] .lut_mask = 64'h9669699696696996;
defparam \o[22] .shared_arith = "off";

dffeas \reg_out[22] (
	.clk(clk),
	.d(\o[22]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[22]~q ),
	.prn(vcc));
defparam \reg_out[22] .is_wysiwyg = "true";
defparam \reg_out[22] .power_up = "low";

cyclonev_lcell_comb \o[14] (
	.dataa(!\reg_out[1]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[14] .extended_lut = "off";
defparam \o[14] .lut_mask = 64'h6996699669966996;
defparam \o[14] .shared_arith = "off";

dffeas \reg_out[14] (
	.clk(clk),
	.d(\o[14]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[14]~q ),
	.prn(vcc));
defparam \reg_out[14] .is_wysiwyg = "true";
defparam \reg_out[14] .power_up = "low";

cyclonev_lcell_comb \o[6] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[5]~q ),
	.datac(!\reg_out[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[6] .extended_lut = "off";
defparam \o[6] .lut_mask = 64'h9696969696969696;
defparam \o[6] .shared_arith = "off";

dffeas \reg_out[6] (
	.clk(clk),
	.d(\o[6]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[6]~q ),
	.prn(vcc));
defparam \reg_out[6] .is_wysiwyg = "true";
defparam \reg_out[6] .power_up = "low";

cyclonev_lcell_comb \o1[0] (
	.dataa(!\reg_out[0]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o1[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o1[0] .extended_lut = "off";
defparam \o1[0] .lut_mask = 64'h6996699669966996;
defparam \o1[0] .shared_arith = "off";

cyclonev_lcell_comb \o[28] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[0]~q ),
	.datac(!\reg_out[5]~q ),
	.datad(!\reg_out[6]~q ),
	.datae(!rd_5_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[28] .extended_lut = "off";
defparam \o[28] .lut_mask = 64'h9669699696696996;
defparam \o[28] .shared_arith = "off";

dffeas \reg_out[28] (
	.clk(clk),
	.d(\o[28]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[28]~q ),
	.prn(vcc));
defparam \reg_out[28] .is_wysiwyg = "true";
defparam \reg_out[28] .power_up = "low";

cyclonev_lcell_comb \o[20] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[7]~q ),
	.datad(!\reg_out[3]~q ),
	.datae(!\reg_out[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[20] .extended_lut = "off";
defparam \o[20] .lut_mask = 64'h9669699696696996;
defparam \o[20] .shared_arith = "off";

dffeas \reg_out[20] (
	.clk(clk),
	.d(\o[20]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[20]~q ),
	.prn(vcc));
defparam \reg_out[20] .is_wysiwyg = "true";
defparam \reg_out[20] .power_up = "low";

cyclonev_lcell_comb \o[12] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[0]~q ),
	.datac(!\reg_out[20]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[12] .extended_lut = "off";
defparam \o[12] .lut_mask = 64'h9696969696969696;
defparam \o[12] .shared_arith = "off";

dffeas \reg_out[12] (
	.clk(clk),
	.d(\o[12]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[12]~q ),
	.prn(vcc));
defparam \reg_out[12] .is_wysiwyg = "true";
defparam \reg_out[12] .power_up = "low";

cyclonev_lcell_comb \o[4] (
	.dataa(!\o1[0]~combout ),
	.datab(!\reg_out[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[4] .extended_lut = "off";
defparam \o[4] .lut_mask = 64'h6666666666666666;
defparam \o[4] .shared_arith = "off";

dffeas \reg_out[4] (
	.clk(clk),
	.d(\o[4]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[4]~q ),
	.prn(vcc));
defparam \reg_out[4] .is_wysiwyg = "true";
defparam \reg_out[4] .power_up = "low";

cyclonev_lcell_comb \o[26] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[1]~q ),
	.datac(!\reg_out[7]~q ),
	.datad(!\o1[0]~combout ),
	.datae(!rd_5_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[26] .extended_lut = "off";
defparam \o[26] .lut_mask = 64'h9669699696696996;
defparam \o[26] .shared_arith = "off";

dffeas \reg_out[26] (
	.clk(clk),
	.d(\o[26]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[26]~q ),
	.prn(vcc));
defparam \reg_out[26] .is_wysiwyg = "true";
defparam \reg_out[26] .power_up = "low";

cyclonev_lcell_comb \o[18]~0 (
	.dataa(!\reg_out[5]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[18]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[18]~0 .extended_lut = "off";
defparam \o[18]~0 .lut_mask = 64'h6996699669966996;
defparam \o[18]~0 .shared_arith = "off";

cyclonev_lcell_comb \o[18] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[0]~q ),
	.datac(!\reg_out[1]~q ),
	.datad(!\o[18]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[18] .extended_lut = "off";
defparam \o[18] .lut_mask = 64'h6996699669966996;
defparam \o[18] .shared_arith = "off";

dffeas \reg_out[18] (
	.clk(clk),
	.d(\o[18]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[18]~q ),
	.prn(vcc));
defparam \reg_out[18] .is_wysiwyg = "true";
defparam \reg_out[18] .power_up = "low";

cyclonev_lcell_comb \o[10] (
	.dataa(!\reg_out[2]~q ),
	.datab(!\reg_out[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[10] .extended_lut = "off";
defparam \o[10] .lut_mask = 64'h6666666666666666;
defparam \o[10] .shared_arith = "off";

dffeas \reg_out[10] (
	.clk(clk),
	.d(\o[10]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[10]~q ),
	.prn(vcc));
defparam \reg_out[10] .is_wysiwyg = "true";
defparam \reg_out[10] .power_up = "low";

cyclonev_lcell_comb \o[2] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[0]~q ),
	.datac(!\reg_out[1]~q ),
	.datad(!\reg_out[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[2] .extended_lut = "off";
defparam \o[2] .lut_mask = 64'h6996699669966996;
defparam \o[2] .shared_arith = "off";

dffeas \reg_out[2] (
	.clk(clk),
	.d(\o[2]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[2]~q ),
	.prn(vcc));
defparam \reg_out[2] .is_wysiwyg = "true";
defparam \reg_out[2] .power_up = "low";

cyclonev_lcell_comb \o[24] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[0]~q ),
	.datac(!\reg_out[5]~q ),
	.datad(!\reg_out[2]~q ),
	.datae(!\reg_out[7]~q ),
	.dataf(!rd_5_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[24] .extended_lut = "off";
defparam \o[24] .lut_mask = 64'h6996966996696996;
defparam \o[24] .shared_arith = "off";

dffeas \reg_out[24] (
	.clk(clk),
	.d(\o[24]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[24]~q ),
	.prn(vcc));
defparam \reg_out[24] .is_wysiwyg = "true";
defparam \reg_out[24] .power_up = "low";

cyclonev_lcell_comb \o[16] (
	.dataa(!\reg_out[4]~q ),
	.datab(!\reg_out[0]~q ),
	.datac(!\reg_out[2]~q ),
	.datad(!\reg_out[3]~q ),
	.datae(!\reg_out[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[16] .extended_lut = "off";
defparam \o[16] .lut_mask = 64'h9669699696696996;
defparam \o[16] .shared_arith = "off";

dffeas \reg_out[16] (
	.clk(clk),
	.d(\o[16]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[16]~q ),
	.prn(vcc));
defparam \reg_out[16] .is_wysiwyg = "true";
defparam \reg_out[16] .power_up = "low";

cyclonev_lcell_comb \o[8] (
	.dataa(!\reg_out[1]~q ),
	.datab(!\reg_out[6]~q ),
	.datac(!\reg_out[7]~q ),
	.datad(!\reg_out[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[8] .extended_lut = "off";
defparam \o[8] .lut_mask = 64'h6996699669966996;
defparam \o[8] .shared_arith = "off";

dffeas \reg_out[8] (
	.clk(clk),
	.d(\o[8]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(sop_4),
	.ena(clk_ena),
	.q(\reg_out[8]~q ),
	.prn(vcc));
defparam \reg_out[8] .is_wysiwyg = "true";
defparam \reg_out[8] .power_up = "low";

cyclonev_lcell_comb \o[0] (
	.dataa(!\reg_out[2]~q ),
	.datab(!\reg_out[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\o[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \o[0] .extended_lut = "off";
defparam \o[0] .lut_mask = 64'h6666666666666666;
defparam \o[0] .shared_arith = "off";

dffeas \reg_out[0] (
	.clk(clk),
	.d(\o[0]~combout ),
	.asdata(vcc),
	.clrn(rst),
	.aload(gnd),
	.sclr(sop_4),
	.sload(gnd),
	.ena(clk_ena),
	.q(\reg_out[0]~q ),
	.prn(vcc));
defparam \reg_out[0] .is_wysiwyg = "true";
defparam \reg_out[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_tx_min_ff (
	q_b_9,
	eop_sft_0,
	q_b_8,
	q_b_4,
	dout_reg_sft_28,
	q_b_0,
	dout_reg_sft_24,
	q_b_5,
	dout_reg_sft_29,
	q_b_1,
	dout_reg_sft_25,
	q_b_6,
	dout_reg_sft_30,
	q_b_2,
	dout_reg_sft_26,
	q_b_7,
	dout_reg_sft_31,
	q_b_3,
	dout_reg_sft_27,
	septy_flag,
	afull_flag,
	aempty_flag,
	altera_tse_reset_synchronizer_chain_out,
	txclk_ena,
	altera_tse_reset_synchronizer_chain_out1,
	tx_empty1,
	tx_data_int_7,
	dreg_1,
	tx_eop_int,
	empty_flag,
	always9,
	col_int,
	always91,
	tx_rden_mii,
	tx_rden_int,
	always92,
	mac_ena,
	sav_flag,
	dreg_11,
	tx_stat_1,
	sop_reg1,
	tx_stat_rden,
	dreg_12,
	tx_stat_0,
	din_s1,
	GND_port,
	clk_32_clk,
	mac_tx_clock_connection_clk,
	mac_misc_connection_ff_tx_crc_fwd)/* synthesis synthesis_greybox=1 */;
output 	q_b_9;
output 	eop_sft_0;
output 	q_b_8;
output 	q_b_4;
output 	dout_reg_sft_28;
output 	q_b_0;
output 	dout_reg_sft_24;
output 	q_b_5;
output 	dout_reg_sft_29;
output 	q_b_1;
output 	dout_reg_sft_25;
output 	q_b_6;
output 	dout_reg_sft_30;
output 	q_b_2;
output 	dout_reg_sft_26;
output 	q_b_7;
output 	dout_reg_sft_31;
output 	q_b_3;
output 	dout_reg_sft_27;
output 	septy_flag;
output 	afull_flag;
output 	aempty_flag;
input 	altera_tse_reset_synchronizer_chain_out;
input 	txclk_ena;
input 	altera_tse_reset_synchronizer_chain_out1;
output 	tx_empty1;
output 	tx_data_int_7;
input 	dreg_1;
output 	tx_eop_int;
output 	empty_flag;
input 	always9;
input 	col_int;
input 	always91;
input 	tx_rden_mii;
input 	tx_rden_int;
input 	always92;
output 	mac_ena;
output 	sav_flag;
input 	dreg_11;
output 	tx_stat_1;
output 	sop_reg1;
input 	tx_stat_rden;
input 	dreg_12;
output 	tx_stat_0;
output 	din_s1;
input 	GND_port;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;
input 	mac_misc_connection_ff_tx_crc_fwd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_RETR|transmit_cnt[0]~q ;
wire \U_RETR|transmit_cnt[1]~q ;
wire \U_RETR|transmit_cnt[2]~q ;
wire \U_RETR|transmit_cnt[3]~q ;
wire \U_RETR|transmit_cnt[4]~q ;
wire \U_RETR|transmit_cnt[5]~q ;
wire \U_RETR|transmit_cnt[6]~q ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ;
wire \TX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[28] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[24] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[29] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[25] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[30] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[26] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[31] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[27] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[20] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[16] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[21] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[17] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[22] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[18] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[23] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[19] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[12] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[8] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[13] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[9] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[14] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[10] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[15] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[11] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[4] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[0] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[5] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[1] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[6] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[2] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[7] ;
wire \TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[3] ;
wire \TX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ;
wire \U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ;
wire \U_RETR|retrans_ena~q ;
wire \U_RETR|buf_wren~q ;
wire \U_RETR|buf_wraddr[0]~q ;
wire \U_RETR|buf_wraddr[1]~q ;
wire \U_RETR|buf_wraddr[2]~q ;
wire \U_RETR|buf_wraddr[3]~q ;
wire \U_RETR|buf_wraddr[4]~q ;
wire \U_RETR|buf_wraddr[5]~q ;
wire \U_RETR|buf_wraddr[6]~q ;
wire \U_RETR|state.STM_TYP_WAIT_COL_1~q ;
wire \U_RETR|state.STM_TYP_RETRANSMIT_SHORT~q ;
wire \U_RETR|Selector4~0_combout ;
wire \U_RETR|short_frm~q ;
wire \U_RETR|Selector1~1_combout ;
wire \U_RETR|Selector5~0_combout ;
wire \U_RETR|always10~0_combout ;
wire \U_RETR|Selector3~0_combout ;
wire \U_RETR|Selector3~2_combout ;
wire \U_RETR|Selector3~3_combout ;
wire \TX_DATA|empty_flag~q ;
wire \always5~0_combout ;
wire \U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_RETR|stat_rden~q ;
wire \comb~0_combout ;
wire \crc_fwd_tmp~q ;
wire \U_SYNC_TX_SHIFT16|std_sync_no_cut|dreg[1]~q ;
wire \TX_DATA|full_flag~q ;
wire \crc_fwd_tmp~0_combout ;
wire \Decoder0~0_combout ;
wire \Decoder0~1_combout ;
wire \Decoder0~2_combout ;
wire \tx_rden~0_combout ;
wire \tx_rden~2_combout ;
wire \tx_rden~1_combout ;
wire \byte_empty~1_combout ;
wire \byte_empty[0]~q ;
wire \byte_empty~0_combout ;
wire \byte_empty[1]~q ;
wire \always4~0_combout ;
wire \eop_sft~1_combout ;
wire \eop_sft~2_combout ;
wire \eop_sft[3]~q ;
wire \always4~2_combout ;
wire \always4~1_combout ;
wire \eop_sft[0]~0_combout ;
wire \eop_sft[2]~q ;
wire \eop_sft[1]~q ;
wire \dout_reg_sft[4]~q ;
wire \dout_reg_sft[12]~q ;
wire \dout_reg_sft[20]~q ;
wire \dout_reg_sft[0]~q ;
wire \dout_reg_sft[8]~q ;
wire \dout_reg_sft[16]~q ;
wire \dout_reg_sft[5]~q ;
wire \dout_reg_sft[13]~q ;
wire \dout_reg_sft[21]~q ;
wire \dout_reg_sft[1]~q ;
wire \dout_reg_sft[9]~q ;
wire \dout_reg_sft[17]~q ;
wire \dout_reg_sft[6]~q ;
wire \dout_reg_sft[14]~q ;
wire \dout_reg_sft[22]~q ;
wire \dout_reg_sft[2]~q ;
wire \dout_reg_sft[10]~q ;
wire \dout_reg_sft[18]~q ;
wire \dout_reg_sft[7]~q ;
wire \dout_reg_sft[15]~q ;
wire \dout_reg_sft[23]~q ;
wire \dout_reg_sft[3]~q ;
wire \dout_reg_sft[11]~q ;
wire \dout_reg_sft[19]~q ;
wire \always6~0_combout ;
wire \sop_reg~1_combout ;
wire \sop_reg~0_combout ;


IoTOctopus_QSYS_altera_tse_a_fifo_13 TX_STATUS(
	.q_b_1(\TX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.q_b_0(\TX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.empty_flag1(empty_flag),
	.comb(\comb~0_combout ),
	.crc_fwd_tmp(\crc_fwd_tmp~q ),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_a_fifo_opt_1246_1 TX_DATA(
	.q_b_34(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.q_b_33(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.q_b_35(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.q_b_32(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.q_b_28(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[28] ),
	.q_b_24(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[24] ),
	.q_b_29(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[29] ),
	.q_b_25(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[25] ),
	.q_b_30(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[30] ),
	.q_b_26(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[26] ),
	.q_b_31(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[31] ),
	.q_b_27(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[27] ),
	.q_b_20(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[20] ),
	.q_b_16(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[16] ),
	.q_b_21(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[21] ),
	.q_b_17(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[17] ),
	.q_b_22(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[22] ),
	.q_b_18(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[18] ),
	.q_b_23(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[23] ),
	.q_b_19(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[19] ),
	.q_b_12(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[12] ),
	.q_b_8(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[8] ),
	.q_b_13(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[13] ),
	.q_b_9(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[9] ),
	.q_b_14(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[14] ),
	.q_b_10(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[10] ),
	.q_b_15(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[15] ),
	.q_b_11(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[11] ),
	.q_b_4(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[4] ),
	.q_b_0(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.q_b_5(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[5] ),
	.q_b_1(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.q_b_6(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[6] ),
	.q_b_2(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.q_b_7(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[7] ),
	.q_b_3(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.septy_flag1(septy_flag),
	.afull_flag1(afull_flag),
	.aempty_flag1(aempty_flag),
	.dreg_1(\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.altera_tse_reset_synchronizer_chain_out1(altera_tse_reset_synchronizer_chain_out1),
	.sav_flag1(sav_flag),
	.empty_flag1(\TX_DATA|empty_flag~q ),
	.always5(\always5~0_combout ),
	.dreg_111(\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_112(\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_113(\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_114(\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_115(\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_116(\U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_117(\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_118(\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_119(\U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_120(\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_121(\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.full_flag1(\TX_DATA|full_flag~q ),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_142 U_SYNC_TX_SHIFT16(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_TX_SHIFT16|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_retransmit_cntl U_RETR(
	.q_b_9(q_b_9),
	.eop_sft_0(eop_sft_0),
	.transmit_cnt_0(\U_RETR|transmit_cnt[0]~q ),
	.transmit_cnt_1(\U_RETR|transmit_cnt[1]~q ),
	.transmit_cnt_2(\U_RETR|transmit_cnt[2]~q ),
	.transmit_cnt_3(\U_RETR|transmit_cnt[3]~q ),
	.transmit_cnt_4(\U_RETR|transmit_cnt[4]~q ),
	.transmit_cnt_5(\U_RETR|transmit_cnt[5]~q ),
	.transmit_cnt_6(\U_RETR|transmit_cnt[6]~q ),
	.clk_ena(txclk_ena),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.retrans_ena1(\U_RETR|retrans_ena~q ),
	.dreg_11(dreg_1),
	.always9(always9),
	.buf_wren1(\U_RETR|buf_wren~q ),
	.buf_wraddr_0(\U_RETR|buf_wraddr[0]~q ),
	.buf_wraddr_1(\U_RETR|buf_wraddr[1]~q ),
	.buf_wraddr_2(\U_RETR|buf_wraddr[2]~q ),
	.buf_wraddr_3(\U_RETR|buf_wraddr[3]~q ),
	.buf_wraddr_4(\U_RETR|buf_wraddr[4]~q ),
	.buf_wraddr_5(\U_RETR|buf_wraddr[5]~q ),
	.buf_wraddr_6(\U_RETR|buf_wraddr[6]~q ),
	.stateSTM_TYP_WAIT_COL_1(\U_RETR|state.STM_TYP_WAIT_COL_1~q ),
	.stateSTM_TYP_RETRANSMIT_SHORT(\U_RETR|state.STM_TYP_RETRANSMIT_SHORT~q ),
	.col_int(col_int),
	.Selector4(\U_RETR|Selector4~0_combout ),
	.short_frm1(\U_RETR|short_frm~q ),
	.always91(always91),
	.tx_rden_mii(tx_rden_mii),
	.Selector1(\U_RETR|Selector1~1_combout ),
	.Selector5(\U_RETR|Selector5~0_combout ),
	.always10(\U_RETR|always10~0_combout ),
	.tx_rden_int(tx_rden_int),
	.Selector3(\U_RETR|Selector3~0_combout ),
	.Selector31(\U_RETR|Selector3~2_combout ),
	.always92(always92),
	.Selector32(\U_RETR|Selector3~3_combout ),
	.mac_ena1(mac_ena),
	.crs(dreg_11),
	.stat_rden1(\U_RETR|stat_rden~q ),
	.tx_stat_rden(tx_stat_rden),
	.GND_port(GND_port),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_141 U_SYNC_HALF_DUPLEX_ENA(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_4 U_RTSM(
	.q_b_9(q_b_9),
	.eop_sft_0(eop_sft_0),
	.transmit_cnt_0(\U_RETR|transmit_cnt[0]~q ),
	.transmit_cnt_1(\U_RETR|transmit_cnt[1]~q ),
	.transmit_cnt_2(\U_RETR|transmit_cnt[2]~q ),
	.transmit_cnt_3(\U_RETR|transmit_cnt[3]~q ),
	.transmit_cnt_4(\U_RETR|transmit_cnt[4]~q ),
	.transmit_cnt_5(\U_RETR|transmit_cnt[5]~q ),
	.transmit_cnt_6(\U_RETR|transmit_cnt[6]~q ),
	.q_b_8(q_b_8),
	.q_b_4(q_b_4),
	.dout_reg_sft_28(dout_reg_sft_28),
	.q_b_0(q_b_0),
	.dout_reg_sft_24(dout_reg_sft_24),
	.q_b_5(q_b_5),
	.dout_reg_sft_29(dout_reg_sft_29),
	.q_b_1(q_b_1),
	.dout_reg_sft_25(dout_reg_sft_25),
	.q_b_6(q_b_6),
	.dout_reg_sft_30(dout_reg_sft_30),
	.q_b_2(q_b_2),
	.dout_reg_sft_26(dout_reg_sft_26),
	.q_b_7(q_b_7),
	.dout_reg_sft_31(dout_reg_sft_31),
	.q_b_3(q_b_3),
	.dout_reg_sft_27(dout_reg_sft_27),
	.buf_wren(\U_RETR|buf_wren~q ),
	.buf_wraddr_0(\U_RETR|buf_wraddr[0]~q ),
	.buf_wraddr_1(\U_RETR|buf_wraddr[1]~q ),
	.buf_wraddr_2(\U_RETR|buf_wraddr[2]~q ),
	.buf_wraddr_3(\U_RETR|buf_wraddr[3]~q ),
	.buf_wraddr_4(\U_RETR|buf_wraddr[4]~q ),
	.buf_wraddr_5(\U_RETR|buf_wraddr[5]~q ),
	.buf_wraddr_6(\U_RETR|buf_wraddr[6]~q ),
	.sop_reg(sop_reg1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_11 U_SYNC_2(
	.dreg_1(\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.din_s1(din_s1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_10 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

cyclonev_lcell_comb \always5~0 (
	.dataa(!\U_RETR|always10~0_combout ),
	.datab(!\tx_rden~0_combout ),
	.datac(!\tx_rden~1_combout ),
	.datad(!\TX_DATA|empty_flag~q ),
	.datae(!\always4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always5~0 .extended_lut = "off";
defparam \always5~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \always5~0 .shared_arith = "off";

cyclonev_lcell_comb \comb~0 (
	.dataa(!empty_flag),
	.datab(!\U_RETR|stat_rden~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \comb~0 .extended_lut = "off";
defparam \comb~0 .lut_mask = 64'h7777777777777777;
defparam \comb~0 .shared_arith = "off";

dffeas crc_fwd_tmp(
	.clk(clk_32_clk),
	.d(\crc_fwd_tmp~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\crc_fwd_tmp~q ),
	.prn(vcc));
defparam crc_fwd_tmp.is_wysiwyg = "true";
defparam crc_fwd_tmp.power_up = "low";

cyclonev_lcell_comb \crc_fwd_tmp~0 (
	.dataa(!\crc_fwd_tmp~q ),
	.datab(!mac_misc_connection_ff_tx_crc_fwd),
	.datac(!dreg_12),
	.datad(!\U_SYNC_TX_SHIFT16|std_sync_no_cut|dreg[1]~q ),
	.datae(!\TX_DATA|full_flag~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\crc_fwd_tmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \crc_fwd_tmp~0 .extended_lut = "off";
defparam \crc_fwd_tmp~0 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \crc_fwd_tmp~0 .shared_arith = "off";

dffeas \eop_sft[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Decoder0~0_combout ),
	.asdata(\eop_sft[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(eop_sft_0),
	.prn(vcc));
defparam \eop_sft[0] .is_wysiwyg = "true";
defparam \eop_sft[0] .power_up = "low";

dffeas \dout_reg_sft[28] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[28] ),
	.asdata(\dout_reg_sft[20]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_28),
	.prn(vcc));
defparam \dout_reg_sft[28] .is_wysiwyg = "true";
defparam \dout_reg_sft[28] .power_up = "low";

dffeas \dout_reg_sft[24] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[24] ),
	.asdata(\dout_reg_sft[16]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_24),
	.prn(vcc));
defparam \dout_reg_sft[24] .is_wysiwyg = "true";
defparam \dout_reg_sft[24] .power_up = "low";

dffeas \dout_reg_sft[29] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[29] ),
	.asdata(\dout_reg_sft[21]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_29),
	.prn(vcc));
defparam \dout_reg_sft[29] .is_wysiwyg = "true";
defparam \dout_reg_sft[29] .power_up = "low";

dffeas \dout_reg_sft[25] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[25] ),
	.asdata(\dout_reg_sft[17]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_25),
	.prn(vcc));
defparam \dout_reg_sft[25] .is_wysiwyg = "true";
defparam \dout_reg_sft[25] .power_up = "low";

dffeas \dout_reg_sft[30] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[30] ),
	.asdata(\dout_reg_sft[22]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_30),
	.prn(vcc));
defparam \dout_reg_sft[30] .is_wysiwyg = "true";
defparam \dout_reg_sft[30] .power_up = "low";

dffeas \dout_reg_sft[26] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[26] ),
	.asdata(\dout_reg_sft[18]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_26),
	.prn(vcc));
defparam \dout_reg_sft[26] .is_wysiwyg = "true";
defparam \dout_reg_sft[26] .power_up = "low";

dffeas \dout_reg_sft[31] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[31] ),
	.asdata(\dout_reg_sft[23]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_31),
	.prn(vcc));
defparam \dout_reg_sft[31] .is_wysiwyg = "true";
defparam \dout_reg_sft[31] .power_up = "low";

dffeas \dout_reg_sft[27] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[27] ),
	.asdata(\dout_reg_sft[19]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(dout_reg_sft_27),
	.prn(vcc));
defparam \dout_reg_sft[27] .is_wysiwyg = "true";
defparam \dout_reg_sft[27] .power_up = "low";

dffeas tx_empty(
	.clk(mac_tx_clock_connection_clk),
	.d(\always6~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_empty1),
	.prn(vcc));
defparam tx_empty.is_wysiwyg = "true";
defparam tx_empty.power_up = "low";

cyclonev_lcell_comb \tx_data_int[7]~0 (
	.dataa(!\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_RETR|retrans_ena~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(tx_data_int_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_data_int[7]~0 .extended_lut = "off";
defparam \tx_data_int[7]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \tx_data_int[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \tx_eop_int~0 (
	.dataa(!q_b_9),
	.datab(!\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_RETR|retrans_ena~q ),
	.datad(!eop_sft_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(tx_eop_int),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_eop_int~0 .extended_lut = "off";
defparam \tx_eop_int~0 .lut_mask = 64'h7DFF7DFF7DFF7DFF;
defparam \tx_eop_int~0 .shared_arith = "off";

dffeas \tx_stat[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_stat_1),
	.prn(vcc));
defparam \tx_stat[1] .is_wysiwyg = "true";
defparam \tx_stat[1] .power_up = "low";

dffeas sop_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(\sop_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sop_reg1),
	.prn(vcc));
defparam sop_reg.is_wysiwyg = "true";
defparam sop_reg.power_up = "low";

dffeas \tx_stat[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_STATUS|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tx_stat_0),
	.prn(vcc));
defparam \tx_stat[0] .is_wysiwyg = "true";
defparam \tx_stat[0] .power_up = "low";

cyclonev_lcell_comb \Decoder0~0 (
	.dataa(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.datab(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~0 .extended_lut = "off";
defparam \Decoder0~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Decoder0~0 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~1 (
	.dataa(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.datab(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~1 .extended_lut = "off";
defparam \Decoder0~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Decoder0~1 .shared_arith = "off";

cyclonev_lcell_comb \Decoder0~2 (
	.dataa(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.datab(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Decoder0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Decoder0~2 .extended_lut = "off";
defparam \Decoder0~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \Decoder0~2 .shared_arith = "off";

cyclonev_lcell_comb \tx_rden~0 (
	.dataa(!txclk_ena),
	.datab(!\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.datac(!dreg_1),
	.datad(!always91),
	.datae(!always9),
	.dataf(!tx_rden_mii),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_rden~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_rden~0 .extended_lut = "off";
defparam \tx_rden~0 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \tx_rden~0 .shared_arith = "off";

cyclonev_lcell_comb \tx_rden~2 (
	.dataa(!txclk_ena),
	.datab(!\U_RETR|short_frm~q ),
	.datac(!\U_RETR|Selector3~0_combout ),
	.datad(!\U_RETR|Selector3~2_combout ),
	.datae(!dreg_1),
	.dataf(!tx_rden_mii),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_rden~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_rden~2 .extended_lut = "off";
defparam \tx_rden~2 .lut_mask = 64'hFFFFFFFFF6F9F9F6;
defparam \tx_rden~2 .shared_arith = "off";

cyclonev_lcell_comb \tx_rden~1 (
	.dataa(!txclk_ena),
	.datab(!\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.datac(!dreg_1),
	.datad(!always91),
	.datae(!always9),
	.dataf(!\tx_rden~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tx_rden~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tx_rden~1 .extended_lut = "off";
defparam \tx_rden~1 .lut_mask = 64'hFFFFFFFFFBFFFFFF;
defparam \tx_rden~1 .shared_arith = "off";

cyclonev_lcell_comb \byte_empty~1 (
	.dataa(!eop_sft_0),
	.datab(!\U_RETR|always10~0_combout ),
	.datac(!\byte_empty[0]~q ),
	.datad(!\tx_rden~0_combout ),
	.datae(!\tx_rden~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_empty~1 .extended_lut = "off";
defparam \byte_empty~1 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \byte_empty~1 .shared_arith = "off";

dffeas \byte_empty[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\byte_empty~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byte_empty[0]~q ),
	.prn(vcc));
defparam \byte_empty[0] .is_wysiwyg = "true";
defparam \byte_empty[0] .power_up = "low";

cyclonev_lcell_comb \byte_empty~0 (
	.dataa(!eop_sft_0),
	.datab(!\U_RETR|always10~0_combout ),
	.datac(!\byte_empty[1]~q ),
	.datad(!\byte_empty[0]~q ),
	.datae(!\tx_rden~0_combout ),
	.dataf(!\tx_rden~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\byte_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \byte_empty~0 .extended_lut = "off";
defparam \byte_empty~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \byte_empty~0 .shared_arith = "off";

dffeas \byte_empty[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\byte_empty~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byte_empty[1]~q ),
	.prn(vcc));
defparam \byte_empty[1] .is_wysiwyg = "true";
defparam \byte_empty[1] .power_up = "low";

cyclonev_lcell_comb \always4~0 (
	.dataa(!\byte_empty[1]~q ),
	.datab(!\byte_empty[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~0 .extended_lut = "off";
defparam \always4~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \always4~0 .shared_arith = "off";

cyclonev_lcell_comb \eop_sft~1 (
	.dataa(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[34] ),
	.datab(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[33] ),
	.datac(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[35] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop_sft~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop_sft~1 .extended_lut = "off";
defparam \eop_sft~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \eop_sft~1 .shared_arith = "off";

cyclonev_lcell_comb \eop_sft~2 (
	.dataa(!\U_RETR|always10~0_combout ),
	.datab(!\tx_rden~0_combout ),
	.datac(!\tx_rden~1_combout ),
	.datad(!\always4~0_combout ),
	.datae(!\eop_sft[3]~q ),
	.dataf(!\eop_sft~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop_sft~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop_sft~2 .extended_lut = "off";
defparam \eop_sft~2 .lut_mask = 64'h96FFFFFFFFFFFFFF;
defparam \eop_sft~2 .shared_arith = "off";

dffeas \eop_sft[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\eop_sft~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\eop_sft[3]~q ),
	.prn(vcc));
defparam \eop_sft[3] .is_wysiwyg = "true";
defparam \eop_sft[3] .power_up = "low";

cyclonev_lcell_comb \always4~2 (
	.dataa(!\U_RETR|Selector4~0_combout ),
	.datab(!txclk_ena),
	.datac(!q_b_9),
	.datad(!\U_RETR|state.STM_TYP_WAIT_COL_1~q ),
	.datae(!\U_RETR|state.STM_TYP_RETRANSMIT_SHORT~q ),
	.dataf(!col_int),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~2 .extended_lut = "off";
defparam \always4~2 .lut_mask = 64'hFFFFFFFBFFFFFFFF;
defparam \always4~2 .shared_arith = "off";

cyclonev_lcell_comb \always4~1 (
	.dataa(!\tx_rden~0_combout ),
	.datab(!\tx_rden~1_combout ),
	.datac(!\always4~0_combout ),
	.datad(!\U_RETR|Selector1~1_combout ),
	.datae(!\U_RETR|Selector5~0_combout ),
	.dataf(!\always4~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always4~1 .extended_lut = "off";
defparam \always4~1 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \always4~1 .shared_arith = "off";

cyclonev_lcell_comb \eop_sft[0]~0 (
	.dataa(!txclk_ena),
	.datab(!\U_SYNC_HALF_DUPLEX_ENA|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_RETR|short_frm~q ),
	.datad(!tx_rden_int),
	.datae(!\U_RETR|always10~0_combout ),
	.dataf(!\U_RETR|Selector3~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\eop_sft[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \eop_sft[0]~0 .extended_lut = "off";
defparam \eop_sft[0]~0 .lut_mask = 64'hFFFFEBFFFFFFBEFF;
defparam \eop_sft[0]~0 .shared_arith = "off";

dffeas \eop_sft[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Decoder0~2_combout ),
	.asdata(\eop_sft[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\eop_sft[2]~q ),
	.prn(vcc));
defparam \eop_sft[2] .is_wysiwyg = "true";
defparam \eop_sft[2] .power_up = "low";

dffeas \eop_sft[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Decoder0~1_combout ),
	.asdata(\eop_sft[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\eop_sft[1]~q ),
	.prn(vcc));
defparam \eop_sft[1] .is_wysiwyg = "true";
defparam \eop_sft[1] .power_up = "low";

dffeas \dout_reg_sft[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[4]~q ),
	.prn(vcc));
defparam \dout_reg_sft[4] .is_wysiwyg = "true";
defparam \dout_reg_sft[4] .power_up = "low";

dffeas \dout_reg_sft[12] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[12] ),
	.asdata(\dout_reg_sft[4]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[12]~q ),
	.prn(vcc));
defparam \dout_reg_sft[12] .is_wysiwyg = "true";
defparam \dout_reg_sft[12] .power_up = "low";

dffeas \dout_reg_sft[20] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[20] ),
	.asdata(\dout_reg_sft[12]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[20]~q ),
	.prn(vcc));
defparam \dout_reg_sft[20] .is_wysiwyg = "true";
defparam \dout_reg_sft[20] .power_up = "low";

dffeas \dout_reg_sft[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[0]~q ),
	.prn(vcc));
defparam \dout_reg_sft[0] .is_wysiwyg = "true";
defparam \dout_reg_sft[0] .power_up = "low";

dffeas \dout_reg_sft[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[8] ),
	.asdata(\dout_reg_sft[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[8]~q ),
	.prn(vcc));
defparam \dout_reg_sft[8] .is_wysiwyg = "true";
defparam \dout_reg_sft[8] .power_up = "low";

dffeas \dout_reg_sft[16] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[16] ),
	.asdata(\dout_reg_sft[8]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[16]~q ),
	.prn(vcc));
defparam \dout_reg_sft[16] .is_wysiwyg = "true";
defparam \dout_reg_sft[16] .power_up = "low";

dffeas \dout_reg_sft[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[5]~q ),
	.prn(vcc));
defparam \dout_reg_sft[5] .is_wysiwyg = "true";
defparam \dout_reg_sft[5] .power_up = "low";

dffeas \dout_reg_sft[13] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[13] ),
	.asdata(\dout_reg_sft[5]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[13]~q ),
	.prn(vcc));
defparam \dout_reg_sft[13] .is_wysiwyg = "true";
defparam \dout_reg_sft[13] .power_up = "low";

dffeas \dout_reg_sft[21] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[21] ),
	.asdata(\dout_reg_sft[13]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[21]~q ),
	.prn(vcc));
defparam \dout_reg_sft[21] .is_wysiwyg = "true";
defparam \dout_reg_sft[21] .power_up = "low";

dffeas \dout_reg_sft[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[1]~q ),
	.prn(vcc));
defparam \dout_reg_sft[1] .is_wysiwyg = "true";
defparam \dout_reg_sft[1] .power_up = "low";

dffeas \dout_reg_sft[9] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[9] ),
	.asdata(\dout_reg_sft[1]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[9]~q ),
	.prn(vcc));
defparam \dout_reg_sft[9] .is_wysiwyg = "true";
defparam \dout_reg_sft[9] .power_up = "low";

dffeas \dout_reg_sft[17] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[17] ),
	.asdata(\dout_reg_sft[9]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[17]~q ),
	.prn(vcc));
defparam \dout_reg_sft[17] .is_wysiwyg = "true";
defparam \dout_reg_sft[17] .power_up = "low";

dffeas \dout_reg_sft[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[6]~q ),
	.prn(vcc));
defparam \dout_reg_sft[6] .is_wysiwyg = "true";
defparam \dout_reg_sft[6] .power_up = "low";

dffeas \dout_reg_sft[14] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[14] ),
	.asdata(\dout_reg_sft[6]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[14]~q ),
	.prn(vcc));
defparam \dout_reg_sft[14] .is_wysiwyg = "true";
defparam \dout_reg_sft[14] .power_up = "low";

dffeas \dout_reg_sft[22] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[22] ),
	.asdata(\dout_reg_sft[14]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[22]~q ),
	.prn(vcc));
defparam \dout_reg_sft[22] .is_wysiwyg = "true";
defparam \dout_reg_sft[22] .power_up = "low";

dffeas \dout_reg_sft[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[2]~q ),
	.prn(vcc));
defparam \dout_reg_sft[2] .is_wysiwyg = "true";
defparam \dout_reg_sft[2] .power_up = "low";

dffeas \dout_reg_sft[10] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[10] ),
	.asdata(\dout_reg_sft[2]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[10]~q ),
	.prn(vcc));
defparam \dout_reg_sft[10] .is_wysiwyg = "true";
defparam \dout_reg_sft[10] .power_up = "low";

dffeas \dout_reg_sft[18] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[18] ),
	.asdata(\dout_reg_sft[10]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[18]~q ),
	.prn(vcc));
defparam \dout_reg_sft[18] .is_wysiwyg = "true";
defparam \dout_reg_sft[18] .power_up = "low";

dffeas \dout_reg_sft[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[7]~q ),
	.prn(vcc));
defparam \dout_reg_sft[7] .is_wysiwyg = "true";
defparam \dout_reg_sft[7] .power_up = "low";

dffeas \dout_reg_sft[15] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[15] ),
	.asdata(\dout_reg_sft[7]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[15]~q ),
	.prn(vcc));
defparam \dout_reg_sft[15] .is_wysiwyg = "true";
defparam \dout_reg_sft[15] .power_up = "low";

dffeas \dout_reg_sft[23] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[23] ),
	.asdata(\dout_reg_sft[15]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[23]~q ),
	.prn(vcc));
defparam \dout_reg_sft[23] .is_wysiwyg = "true";
defparam \dout_reg_sft[23] .power_up = "low";

dffeas \dout_reg_sft[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always4~1_combout ),
	.q(\dout_reg_sft[3]~q ),
	.prn(vcc));
defparam \dout_reg_sft[3] .is_wysiwyg = "true";
defparam \dout_reg_sft[3] .power_up = "low";

dffeas \dout_reg_sft[11] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[11] ),
	.asdata(\dout_reg_sft[3]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[11]~q ),
	.prn(vcc));
defparam \dout_reg_sft[11] .is_wysiwyg = "true";
defparam \dout_reg_sft[11] .power_up = "low";

dffeas \dout_reg_sft[19] (
	.clk(mac_tx_clock_connection_clk),
	.d(\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[19] ),
	.asdata(\dout_reg_sft[11]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\always4~1_combout ),
	.ena(\eop_sft[0]~0_combout ),
	.q(\dout_reg_sft[19]~q ),
	.prn(vcc));
defparam \dout_reg_sft[19] .is_wysiwyg = "true";
defparam \dout_reg_sft[19] .power_up = "low";

cyclonev_lcell_comb \always6~0 (
	.dataa(!aempty_flag),
	.datab(!empty_flag),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always6~0 .extended_lut = "off";
defparam \always6~0 .lut_mask = 64'h7777777777777777;
defparam \always6~0 .shared_arith = "off";

cyclonev_lcell_comb \sop_reg~1 (
	.dataa(!\TX_DATA|empty_flag~q ),
	.datab(!\always4~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_reg~1 .extended_lut = "off";
defparam \sop_reg~1 .lut_mask = 64'h7777777777777777;
defparam \sop_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \sop_reg~0 (
	.dataa(!\U_RETR|always10~0_combout ),
	.datab(!\tx_rden~0_combout ),
	.datac(!\tx_rden~1_combout ),
	.datad(!sop_reg1),
	.datae(!\TX_DATA|U_RAM|altsyncram_component|auto_generated|q_b[32] ),
	.dataf(!\sop_reg~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sop_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sop_reg~0 .extended_lut = "off";
defparam \sop_reg~0 .lut_mask = 64'h96FFFFFFFFFFFFFF;
defparam \sop_reg~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_141 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_141 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_141 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_142 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_142 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_142 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_10 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_144 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_153 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_152 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_151 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_150 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_149 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_148 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_147 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_146 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_145 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_143 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_143 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_143 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_143 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_144 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_144 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_144 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_145 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_145 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_145 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_146 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_146 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_146 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_147 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_147 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_147 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_148 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_148 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_148 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_149 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_149 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_149 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_150 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_150 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_150 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_151 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_151 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_151 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_152 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_152 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_152 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_153 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_153 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_153 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_11 (
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	altera_tse_reset_synchronizer_chain_out,
	din_s1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	altera_tse_reset_synchronizer_chain_out;
output 	din_s1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_155 \sync[10].u (
	.dreg_1(dreg_1),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.din_s1(din_s1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_164 \sync[9].u (
	.dreg_1(dreg_110),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_163 \sync[8].u (
	.dreg_1(dreg_19),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_162 \sync[7].u (
	.dreg_1(dreg_18),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_161 \sync[6].u (
	.dreg_1(dreg_17),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_160 \sync[5].u (
	.dreg_1(dreg_16),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_159 \sync[4].u (
	.dreg_1(dreg_15),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_158 \sync[3].u (
	.dreg_1(dreg_14),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_157 \sync[2].u (
	.dreg_1(dreg_13),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_156 \sync[1].u (
	.dreg_1(dreg_12),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_154 \sync[0].u (
	.dreg_1(dreg_11),
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_154 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_154 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_154 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_155 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	din_s1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
output 	din_s1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_155 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.din_s11(din_s1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_155 (
	dreg_1,
	reset_n,
	din_s11,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
output 	din_s11;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(din_s11),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(din_s11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_156 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_156 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_156 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_157 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_157 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_157 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_158 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_158 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_158 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_159 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_159 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_159 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_160 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_160 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_160 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_161 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_161 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_161 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_162 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_162 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_162 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_163 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_163 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_163 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_164 (
	dreg_1,
	altera_tse_reset_synchronizer_chain_out,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	altera_tse_reset_synchronizer_chain_out;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_164 std_sync_no_cut(
	.dreg_1(dreg_1),
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_164 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_a_fifo_13 (
	q_b_1,
	q_b_0,
	altera_tse_reset_synchronizer_chain_out,
	altera_tse_reset_synchronizer_chain_out1,
	empty_flag1,
	comb,
	crc_fwd_tmp,
	GND_port,
	clk_32_clk,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
input 	altera_tse_reset_synchronizer_chain_out;
input 	altera_tse_reset_synchronizer_chain_out1;
output 	empty_flag1;
input 	comb;
input 	crc_fwd_tmp;
input 	GND_port;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_RD|b_out[3]~q ;
wire \U_RD|b_out[4]~q ;
wire \U_RD|b_out[1]~q ;
wire \U_RD|b_out[2]~q ;
wire \U_RD|b_out[0]~q ;
wire \U_RD|b_out[5]~q ;
wire \U_RD|b_out[6]~q ;
wire \U_RD|b_out[7]~q ;
wire \U_RD|b_out[8]~q ;
wire \U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_WRT|b_out[0]~q ;
wire \U_WRT|b_out[1]~q ;
wire \U_WRT|b_out[2]~q ;
wire \U_WRT|b_out[3]~q ;
wire \U_WRT|b_out[4]~q ;
wire \U_WRT|b_out[5]~q ;
wire \U_WRT|b_out[6]~q ;
wire \U_WRT|b_out[7]~q ;
wire \U_WRT|b_out[8]~q ;
wire \U_WRT|g_out[3]~q ;
wire \U_WRT|g_out[4]~q ;
wire \U_WRT|g_out[5]~q ;
wire \U_WRT|g_out[6]~q ;
wire \U_WRT|g_out[7]~q ;
wire \U_WRT|g_out[8]~q ;
wire \U_WRT|g_out[1]~q ;
wire \U_WRT|g_out[2]~q ;
wire \U_WRT|g_out[0]~q ;
wire \ff_wr_binval[7]~0_combout ;
wire \ff_wr_binval[5]~1_combout ;
wire \ff_wr_binval[5]~3_combout ;
wire \ff_wr_binval[3]~4_combout ;
wire \wr_b_rptr[4]~q ;
wire \ff_wr_binval[3]~2_combout ;
wire \wr_b_rptr[3]~q ;
wire \ff_wr_binval[1]~6_combout ;
wire \wr_b_rptr[2]~q ;
wire \ff_wr_binval[0]~5_combout ;
wire \wr_b_rptr[1]~q ;
wire \ff_wr_binval[0]~combout ;
wire \wr_b_rptr[0]~q ;
wire \ptr_rck_diff[0]~18 ;
wire \ptr_rck_diff[0]~19 ;
wire \ptr_rck_diff[1]~10 ;
wire \ptr_rck_diff[1]~11 ;
wire \ptr_rck_diff[2]~14 ;
wire \ptr_rck_diff[2]~15 ;
wire \ptr_rck_diff[3]~2 ;
wire \ptr_rck_diff[3]~3 ;
wire \ptr_rck_diff[4]~5_sumout ;
wire \wr_b_rptr[5]~q ;
wire \ptr_rck_diff[4]~6 ;
wire \ptr_rck_diff[4]~7 ;
wire \ptr_rck_diff[5]~21_sumout ;
wire \wr_b_rptr[6]~q ;
wire \ptr_rck_diff[5]~22 ;
wire \ptr_rck_diff[5]~23 ;
wire \ptr_rck_diff[6]~25_sumout ;
wire \wr_b_rptr[7]~q ;
wire \ptr_rck_diff[6]~26 ;
wire \ptr_rck_diff[6]~27 ;
wire \ptr_rck_diff[7]~29_sumout ;
wire \wr_b_rptr[8]~q ;
wire \ptr_rck_diff[7]~30 ;
wire \ptr_rck_diff[7]~31 ;
wire \ptr_rck_diff[8]~33_sumout ;
wire \ptr_rck_diff[3]~1_sumout ;
wire \ptr_rck_diff[1]~9_sumout ;
wire \ptr_rck_diff[2]~13_sumout ;
wire \rden_reg~q ;
wire \ptr_rck_diff[0]~17_sumout ;
wire \empty_flag~1_combout ;
wire \empty_flag~0_combout ;


IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_2 U_RAM(
	.q_b_1(q_b_1),
	.q_b_0(q_b_0),
	.b_out_3(\U_RD|b_out[3]~q ),
	.b_out_4(\U_RD|b_out[4]~q ),
	.b_out_1(\U_RD|b_out[1]~q ),
	.b_out_2(\U_RD|b_out[2]~q ),
	.b_out_0(\U_RD|b_out[0]~q ),
	.b_out_5(\U_RD|b_out[5]~q ),
	.b_out_6(\U_RD|b_out[6]~q ),
	.b_out_7(\U_RD|b_out[7]~q ),
	.b_out_8(\U_RD|b_out[8]~q ),
	.crc_fwd_tmp(crc_fwd_tmp),
	.b_out_01(\U_WRT|b_out[0]~q ),
	.b_out_11(\U_WRT|b_out[1]~q ),
	.b_out_21(\U_WRT|b_out[2]~q ),
	.b_out_31(\U_WRT|b_out[3]~q ),
	.b_out_41(\U_WRT|b_out[4]~q ),
	.b_out_51(\U_WRT|b_out[5]~q ),
	.b_out_61(\U_WRT|b_out[6]~q ),
	.b_out_71(\U_WRT|b_out[7]~q ),
	.b_out_81(\U_WRT|b_out[8]~q ),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_13 U_SYNC_2(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_5 U_RD(
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.b_out_3(\U_RD|b_out[3]~q ),
	.b_out_4(\U_RD|b_out[4]~q ),
	.b_out_1(\U_RD|b_out[1]~q ),
	.b_out_2(\U_RD|b_out[2]~q ),
	.comb(comb),
	.b_out_0(\U_RD|b_out[0]~q ),
	.b_out_5(\U_RD|b_out[5]~q ),
	.b_out_6(\U_RD|b_out[6]~q ),
	.b_out_7(\U_RD|b_out[7]~q ),
	.b_out_8(\U_RD|b_out[8]~q ),
	.clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_6 U_WRT(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ));

dffeas empty_flag(
	.clk(mac_tx_clock_connection_clk),
	.d(\empty_flag~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_flag1),
	.prn(vcc));
defparam empty_flag.is_wysiwyg = "true";
defparam empty_flag.power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[7]~0 (
	.dataa(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[7]~0 .extended_lut = "off";
defparam \ff_wr_binval[7]~0 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \ff_wr_binval[5]~1 (
	.dataa(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\ff_wr_binval[7]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[5]~1 .extended_lut = "off";
defparam \ff_wr_binval[5]~1 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \ff_wr_binval[5]~3 (
	.dataa(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\ff_wr_binval[5]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[5]~3 .extended_lut = "off";
defparam \ff_wr_binval[5]~3 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \ff_wr_binval[3]~4 (
	.dataa(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\ff_wr_binval[5]~3_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~4 .extended_lut = "off";
defparam \ff_wr_binval[3]~4 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[3]~4 .shared_arith = "off";

dffeas \wr_b_rptr[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[3]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[4]~q ),
	.prn(vcc));
defparam \wr_b_rptr[4] .is_wysiwyg = "true";
defparam \wr_b_rptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[3]~2 (
	.dataa(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\ff_wr_binval[5]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~2 .extended_lut = "off";
defparam \ff_wr_binval[3]~2 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[3]~2 .shared_arith = "off";

dffeas \wr_b_rptr[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[3]~q ),
	.prn(vcc));
defparam \wr_b_rptr[3] .is_wysiwyg = "true";
defparam \wr_b_rptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[1]~6 (
	.dataa(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\ff_wr_binval[3]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[1]~6 .extended_lut = "off";
defparam \ff_wr_binval[1]~6 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[1]~6 .shared_arith = "off";

dffeas \wr_b_rptr[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[1]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[2]~q ),
	.prn(vcc));
defparam \wr_b_rptr[2] .is_wysiwyg = "true";
defparam \wr_b_rptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0]~5 (
	.dataa(!\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ff_wr_binval[3]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0]~5 .extended_lut = "off";
defparam \ff_wr_binval[0]~5 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[0]~5 .shared_arith = "off";

dffeas \wr_b_rptr[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[0]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[1]~q ),
	.prn(vcc));
defparam \wr_b_rptr[1] .is_wysiwyg = "true";
defparam \wr_b_rptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0] (
	.dataa(!\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ff_wr_binval[3]~2_combout ),
	.datad(!\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0] .extended_lut = "off";
defparam \ff_wr_binval[0] .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[0] .shared_arith = "off";

dffeas \wr_b_rptr[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[0]~q ),
	.prn(vcc));
defparam \wr_b_rptr[0] .is_wysiwyg = "true";
defparam \wr_b_rptr[0] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[0]~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[0]~q ),
	.datad(!\U_RD|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\ptr_rck_diff[0]~17_sumout ),
	.cout(\ptr_rck_diff[0]~18 ),
	.shareout(\ptr_rck_diff[0]~19 ));
defparam \ptr_rck_diff[0]~17 .extended_lut = "off";
defparam \ptr_rck_diff[0]~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[0]~17 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[1]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[1]~q ),
	.datad(!\U_RD|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[0]~18 ),
	.sharein(\ptr_rck_diff[0]~19 ),
	.combout(),
	.sumout(\ptr_rck_diff[1]~9_sumout ),
	.cout(\ptr_rck_diff[1]~10 ),
	.shareout(\ptr_rck_diff[1]~11 ));
defparam \ptr_rck_diff[1]~9 .extended_lut = "off";
defparam \ptr_rck_diff[1]~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[1]~9 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[2]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[2]~q ),
	.datad(!\U_RD|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[1]~10 ),
	.sharein(\ptr_rck_diff[1]~11 ),
	.combout(),
	.sumout(\ptr_rck_diff[2]~13_sumout ),
	.cout(\ptr_rck_diff[2]~14 ),
	.shareout(\ptr_rck_diff[2]~15 ));
defparam \ptr_rck_diff[2]~13 .extended_lut = "off";
defparam \ptr_rck_diff[2]~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[2]~13 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[3]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[3]~q ),
	.datad(!\U_RD|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[2]~14 ),
	.sharein(\ptr_rck_diff[2]~15 ),
	.combout(),
	.sumout(\ptr_rck_diff[3]~1_sumout ),
	.cout(\ptr_rck_diff[3]~2 ),
	.shareout(\ptr_rck_diff[3]~3 ));
defparam \ptr_rck_diff[3]~1 .extended_lut = "off";
defparam \ptr_rck_diff[3]~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[3]~1 .shared_arith = "on";

cyclonev_lcell_comb \ptr_rck_diff[4]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[4]~q ),
	.datad(!\U_RD|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[3]~2 ),
	.sharein(\ptr_rck_diff[3]~3 ),
	.combout(),
	.sumout(\ptr_rck_diff[4]~5_sumout ),
	.cout(\ptr_rck_diff[4]~6 ),
	.shareout(\ptr_rck_diff[4]~7 ));
defparam \ptr_rck_diff[4]~5 .extended_lut = "off";
defparam \ptr_rck_diff[4]~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[4]~5 .shared_arith = "on";

dffeas \wr_b_rptr[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[5]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[5]~q ),
	.prn(vcc));
defparam \wr_b_rptr[5] .is_wysiwyg = "true";
defparam \wr_b_rptr[5] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[5]~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[5]~q ),
	.datad(!\U_RD|b_out[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[4]~6 ),
	.sharein(\ptr_rck_diff[4]~7 ),
	.combout(),
	.sumout(\ptr_rck_diff[5]~21_sumout ),
	.cout(\ptr_rck_diff[5]~22 ),
	.shareout(\ptr_rck_diff[5]~23 ));
defparam \ptr_rck_diff[5]~21 .extended_lut = "off";
defparam \ptr_rck_diff[5]~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[5]~21 .shared_arith = "on";

dffeas \wr_b_rptr[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[5]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[6]~q ),
	.prn(vcc));
defparam \wr_b_rptr[6] .is_wysiwyg = "true";
defparam \wr_b_rptr[6] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[6]~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[6]~q ),
	.datad(!\U_RD|b_out[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[5]~22 ),
	.sharein(\ptr_rck_diff[5]~23 ),
	.combout(),
	.sumout(\ptr_rck_diff[6]~25_sumout ),
	.cout(\ptr_rck_diff[6]~26 ),
	.shareout(\ptr_rck_diff[6]~27 ));
defparam \ptr_rck_diff[6]~25 .extended_lut = "off";
defparam \ptr_rck_diff[6]~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[6]~25 .shared_arith = "on";

dffeas \wr_b_rptr[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[7]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[7]~q ),
	.prn(vcc));
defparam \wr_b_rptr[7] .is_wysiwyg = "true";
defparam \wr_b_rptr[7] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[7]~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[7]~q ),
	.datad(!\U_RD|b_out[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[6]~26 ),
	.sharein(\ptr_rck_diff[6]~27 ),
	.combout(),
	.sumout(\ptr_rck_diff[7]~29_sumout ),
	.cout(\ptr_rck_diff[7]~30 ),
	.shareout(\ptr_rck_diff[7]~31 ));
defparam \ptr_rck_diff[7]~29 .extended_lut = "off";
defparam \ptr_rck_diff[7]~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \ptr_rck_diff[7]~29 .shared_arith = "on";

dffeas \wr_b_rptr[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[8]~q ),
	.prn(vcc));
defparam \wr_b_rptr[8] .is_wysiwyg = "true";
defparam \wr_b_rptr[8] .power_up = "low";

cyclonev_lcell_comb \ptr_rck_diff[8]~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[8]~q ),
	.datad(!\U_RD|b_out[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\ptr_rck_diff[7]~30 ),
	.sharein(\ptr_rck_diff[7]~31 ),
	.combout(),
	.sumout(\ptr_rck_diff[8]~33_sumout ),
	.cout(),
	.shareout());
defparam \ptr_rck_diff[8]~33 .extended_lut = "off";
defparam \ptr_rck_diff[8]~33 .lut_mask = 64'h0000000000000FF0;
defparam \ptr_rck_diff[8]~33 .shared_arith = "on";

dffeas rden_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(comb),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rden_reg~q ),
	.prn(vcc));
defparam rden_reg.is_wysiwyg = "true";
defparam rden_reg.power_up = "low";

cyclonev_lcell_comb \empty_flag~1 (
	.dataa(!\ptr_rck_diff[3]~1_sumout ),
	.datab(!\ptr_rck_diff[1]~9_sumout ),
	.datac(!\ptr_rck_diff[2]~13_sumout ),
	.datad(!\rden_reg~q ),
	.datae(!\ptr_rck_diff[0]~17_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~1 .extended_lut = "off";
defparam \empty_flag~1 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \empty_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \empty_flag~0 (
	.dataa(!\ptr_rck_diff[4]~5_sumout ),
	.datab(!\ptr_rck_diff[5]~21_sumout ),
	.datac(!\ptr_rck_diff[6]~25_sumout ),
	.datad(!\ptr_rck_diff[7]~29_sumout ),
	.datae(!\ptr_rck_diff[8]~33_sumout ),
	.dataf(!\empty_flag~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~0 .extended_lut = "off";
defparam \empty_flag~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \empty_flag~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_13 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	g_out_3,
	g_out_4,
	g_out_5,
	g_out_6,
	g_out_7,
	g_out_8,
	g_out_1,
	g_out_2,
	g_out_0,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
input 	g_out_3;
input 	g_out_4;
input 	g_out_5;
input 	g_out_6;
input 	g_out_7;
input 	g_out_8;
input 	g_out_1;
input 	g_out_2;
input 	g_out_0;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_182 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.g_out_8(g_out_8),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_181 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.g_out_7(g_out_7),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_175 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.g_out_1(g_out_1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_174 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.g_out_0(g_out_0),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_180 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.g_out_6(g_out_6),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_179 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.g_out_5(g_out_5),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_178 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.g_out_4(g_out_4),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_177 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.g_out_3(g_out_3),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_176 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.g_out_2(g_out_2),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_174 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_0,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_0;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_174 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_0),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_174 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_175 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_175 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_175 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_176 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_2,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_2;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_176 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_2),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_176 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_177 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_3,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_3;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_177 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_3),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_177 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_178 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_4,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_4;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_178 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_4),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_178 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_179 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_5,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_5;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_179 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_5),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_179 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_180 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_6,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_6;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_180 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_6),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_180 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_181 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_7,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_7;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_181 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_7),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_181 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_182 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_8,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_8;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_182 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_8),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_182 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_2 (
	q_b_1,
	q_b_0,
	b_out_3,
	b_out_4,
	b_out_1,
	b_out_2,
	b_out_0,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	crc_fwd_tmp,
	b_out_01,
	b_out_11,
	b_out_21,
	b_out_31,
	b_out_41,
	b_out_51,
	b_out_61,
	b_out_71,
	b_out_81,
	GND_port,
	clk_32_clk,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
input 	b_out_3;
input 	b_out_4;
input 	b_out_1;
input 	b_out_2;
input 	b_out_0;
input 	b_out_5;
input 	b_out_6;
input 	b_out_7;
input 	b_out_8;
input 	crc_fwd_tmp;
input 	b_out_01;
input 	b_out_11;
input 	b_out_21;
input 	b_out_31;
input 	b_out_41;
input 	b_out_51;
input 	b_out_61;
input 	b_out_71;
input 	b_out_81;
input 	GND_port;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_4 altsyncram_component(
	.q_b({q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_unconnected_wire_35,q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,
q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,
q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,
q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_1,q_b_0}),
	.address_b({gnd,gnd,b_out_8,b_out_7,b_out_6,b_out_5,b_out_4,b_out_3,b_out_2,b_out_1,b_out_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,crc_fwd_tmp,GND_port}),
	.address_a({gnd,gnd,b_out_81,b_out_71,b_out_61,b_out_51,b_out_41,b_out_31,b_out_21,b_out_11,b_out_01}),
	.clock0(clk_32_clk),
	.clock1(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altsyncram_4 (
	q_b,
	address_b,
	data_a,
	address_a,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	[10:0] address_b;
input 	[39:0] data_a;
input 	[10:0] address_a;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_n0o1 auto_generated(
	.q_b({q_b[1],q_b[0]}),
	.address_b({address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[1],data_a[0]}),
	.address_a({address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0),
	.clock1(clock1));

endmodule

module IoTOctopus_QSYS_altsyncram_n0o1 (
	q_b,
	address_b,
	data_a,
	address_a,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[1:0] q_b;
input 	[8:0] address_b;
input 	[1:0] data_a;
input 	[8:0] address_a;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a1(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_13:TX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_n0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 9;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 511;
defparam ram_block1a1.port_a_logical_ram_depth = 512;
defparam ram_block1a1.port_a_logical_ram_width = 2;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 9;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 511;
defparam ram_block1a1.port_b_logical_ram_depth = 512;
defparam ram_block1a1.port_b_logical_ram_width = 2;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_13:TX_STATUS|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_n0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 9;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 511;
defparam ram_block1a0.port_a_logical_ram_depth = 512;
defparam ram_block1a0.port_a_logical_ram_width = 2;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 9;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 511;
defparam ram_block1a0.port_b_logical_ram_depth = 512;
defparam ram_block1a0.port_b_logical_ram_width = 2;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_5 (
	reset,
	b_out_3,
	b_out_4,
	b_out_1,
	b_out_2,
	comb,
	b_out_0,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	b_out_3;
output 	b_out_4;
output 	b_out_1;
output 	b_out_2;
input 	comb;
output 	b_out_0;
output 	b_out_5;
output 	b_out_6;
output 	b_out_7;
output 	b_out_8;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~17_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \b_int[4]~q ;
wire \Add0~6 ;
wire \Add0~21_sumout ;
wire \b_int[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \b_int[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \b_int[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \b_int[8]~q ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \b_int~0_combout ;
wire \b_int[0]~q ;
wire \Add0~18 ;
wire \Add0~9_sumout ;
wire \b_int[1]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \b_int[2]~q ;
wire \Add0~14 ;
wire \Add0~1_sumout ;
wire \b_int[3]~q ;
wire \b_out[0]~0_combout ;


dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[5] (
	.clk(clk),
	.d(\b_int[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[6] (
	.clk(clk),
	.d(\b_int[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[7] (
	.clk(clk),
	.d(\b_int[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \b_int[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[5]~q ),
	.prn(vcc));
defparam \b_int[5] .is_wysiwyg = "true";
defparam \b_int[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \b_int[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[6]~q ),
	.prn(vcc));
defparam \b_int[6] .is_wysiwyg = "true";
defparam \b_int[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \b_int[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[7]~q ),
	.prn(vcc));
defparam \b_int[7] .is_wysiwyg = "true";
defparam \b_int[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \b_int[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[8]~q ),
	.prn(vcc));
defparam \b_int[8] .is_wysiwyg = "true";
defparam \b_int[8] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[2]~q ),
	.datac(!\b_int[3]~q ),
	.datad(!\b_int[7]~q ),
	.datae(!\b_int[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\b_int[4]~q ),
	.datab(!\b_int[5]~q ),
	.datac(!\b_int[6]~q ),
	.datad(!\b_int[8]~q ),
	.datae(!\LessThan0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \b_int~0 (
	.dataa(!\Add0~17_sumout ),
	.datab(!\LessThan0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int~0 .extended_lut = "off";
defparam \b_int~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \b_int~0 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

dffeas \b_int[3] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~1_combout ),
	.sload(gnd),
	.ena(comb),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_6 (
	altera_tse_reset_synchronizer_chain_out,
	b_out_0,
	b_out_1,
	b_out_2,
	b_out_3,
	b_out_4,
	b_out_5,
	b_out_6,
	b_out_7,
	b_out_8,
	g_out_3,
	g_out_4,
	g_out_5,
	g_out_6,
	g_out_7,
	g_out_8,
	g_out_1,
	g_out_2,
	g_out_0)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	b_out_0;
output 	b_out_1;
output 	b_out_2;
output 	b_out_3;
output 	b_out_4;
output 	b_out_5;
output 	b_out_6;
output 	b_out_7;
output 	b_out_8;
output 	g_out_3;
output 	g_out_4;
output 	g_out_5;
output 	g_out_6;
output 	g_out_7;
output 	g_out_8;
output 	g_out_1;
output 	g_out_2;
output 	g_out_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \b_out[1]~0_combout ;
wire \b_out[2]~1_combout ;
wire \b_out[3]~2_combout ;
wire \b_out[4]~3_combout ;
wire \b_out[5]~4_combout ;
wire \b_out[6]~5_combout ;
wire \b_out[7]~6_combout ;
wire \b_out[8]~7_combout ;
wire \g_out[3]~0_combout ;
wire \g_out[4]~1_combout ;
wire \g_out[5]~2_combout ;
wire \g_out[6]~3_combout ;
wire \g_out[7]~4_combout ;
wire \g_out[8]~5_combout ;
wire \g_out[1]~6_combout ;
wire \g_out[2]~7_combout ;


dffeas \b_out[0] (
	.clk(gnd),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[1] (
	.clk(gnd),
	.d(\b_out[1]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[2] (
	.clk(gnd),
	.d(\b_out[2]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[3] (
	.clk(gnd),
	.d(\b_out[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[4] (
	.clk(gnd),
	.d(\b_out[4]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[5] (
	.clk(gnd),
	.d(\b_out[5]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[6] (
	.clk(gnd),
	.d(\b_out[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[7] (
	.clk(gnd),
	.d(\b_out[7]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[8] (
	.clk(gnd),
	.d(\b_out[8]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

dffeas \g_out[3] (
	.clk(gnd),
	.d(\g_out[3]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[4] (
	.clk(gnd),
	.d(\g_out[4]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[5] (
	.clk(gnd),
	.d(\g_out[5]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_5),
	.prn(vcc));
defparam \g_out[5] .is_wysiwyg = "true";
defparam \g_out[5] .power_up = "low";

dffeas \g_out[6] (
	.clk(gnd),
	.d(\g_out[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_6),
	.prn(vcc));
defparam \g_out[6] .is_wysiwyg = "true";
defparam \g_out[6] .power_up = "low";

dffeas \g_out[7] (
	.clk(gnd),
	.d(\g_out[7]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_7),
	.prn(vcc));
defparam \g_out[7] .is_wysiwyg = "true";
defparam \g_out[7] .power_up = "low";

dffeas \g_out[8] (
	.clk(gnd),
	.d(\g_out[8]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_8),
	.prn(vcc));
defparam \g_out[8] .is_wysiwyg = "true";
defparam \g_out[8] .power_up = "low";

dffeas \g_out[1] (
	.clk(gnd),
	.d(\g_out[1]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[2] (
	.clk(gnd),
	.d(\g_out[2]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[0] (
	.clk(gnd),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

cyclonev_lcell_comb \b_out[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[1]~0 .extended_lut = "off";
defparam \b_out[1]~0 .lut_mask = 64'h0000000000000000;
defparam \b_out[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \b_out[2]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[2]~1 .extended_lut = "off";
defparam \b_out[2]~1 .lut_mask = 64'h0000000000000000;
defparam \b_out[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \b_out[3]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[3]~2 .extended_lut = "off";
defparam \b_out[3]~2 .lut_mask = 64'h0000000000000000;
defparam \b_out[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \b_out[4]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[4]~3 .extended_lut = "off";
defparam \b_out[4]~3 .lut_mask = 64'h0000000000000000;
defparam \b_out[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \b_out[5]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[5]~4 .extended_lut = "off";
defparam \b_out[5]~4 .lut_mask = 64'h0000000000000000;
defparam \b_out[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \b_out[6]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[6]~5 .extended_lut = "off";
defparam \b_out[6]~5 .lut_mask = 64'h0000000000000000;
defparam \b_out[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \b_out[7]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[7]~6 .extended_lut = "off";
defparam \b_out[7]~6 .lut_mask = 64'h0000000000000000;
defparam \b_out[7]~6 .shared_arith = "off";

cyclonev_lcell_comb \b_out[8]~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[8]~7 .extended_lut = "off";
defparam \b_out[8]~7 .lut_mask = 64'h0000000000000000;
defparam \b_out[8]~7 .shared_arith = "off";

cyclonev_lcell_comb \g_out[3]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[3]~0 .extended_lut = "off";
defparam \g_out[3]~0 .lut_mask = 64'h0000000000000000;
defparam \g_out[3]~0 .shared_arith = "off";

cyclonev_lcell_comb \g_out[4]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[4]~1 .extended_lut = "off";
defparam \g_out[4]~1 .lut_mask = 64'h0000000000000000;
defparam \g_out[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \g_out[5]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[5]~2 .extended_lut = "off";
defparam \g_out[5]~2 .lut_mask = 64'h0000000000000000;
defparam \g_out[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \g_out[6]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[6]~3 .extended_lut = "off";
defparam \g_out[6]~3 .lut_mask = 64'h0000000000000000;
defparam \g_out[6]~3 .shared_arith = "off";

cyclonev_lcell_comb \g_out[7]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[7]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[7]~4 .extended_lut = "off";
defparam \g_out[7]~4 .lut_mask = 64'h0000000000000000;
defparam \g_out[7]~4 .shared_arith = "off";

cyclonev_lcell_comb \g_out[8]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[8]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[8]~5 .extended_lut = "off";
defparam \g_out[8]~5 .lut_mask = 64'h0000000000000000;
defparam \g_out[8]~5 .shared_arith = "off";

cyclonev_lcell_comb \g_out[1]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[1]~6 .extended_lut = "off";
defparam \g_out[1]~6 .lut_mask = 64'h0000000000000000;
defparam \g_out[1]~6 .shared_arith = "off";

cyclonev_lcell_comb \g_out[2]~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[2]~7 .extended_lut = "off";
defparam \g_out[2]~7 .lut_mask = 64'h0000000000000000;
defparam \g_out[2]~7 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_a_fifo_opt_1246_1 (
	q_b_34,
	q_b_33,
	q_b_35,
	q_b_32,
	q_b_28,
	q_b_24,
	q_b_29,
	q_b_25,
	q_b_30,
	q_b_26,
	q_b_31,
	q_b_27,
	q_b_20,
	q_b_16,
	q_b_21,
	q_b_17,
	q_b_22,
	q_b_18,
	q_b_23,
	q_b_19,
	q_b_12,
	q_b_8,
	q_b_13,
	q_b_9,
	q_b_14,
	q_b_10,
	q_b_15,
	q_b_11,
	q_b_4,
	q_b_0,
	q_b_5,
	q_b_1,
	q_b_6,
	q_b_2,
	q_b_7,
	q_b_3,
	septy_flag1,
	afull_flag1,
	aempty_flag1,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	altera_tse_reset_synchronizer_chain_out,
	altera_tse_reset_synchronizer_chain_out1,
	sav_flag1,
	empty_flag1,
	always5,
	dreg_111,
	dreg_112,
	dreg_113,
	dreg_114,
	dreg_115,
	dreg_116,
	dreg_117,
	dreg_118,
	dreg_119,
	dreg_120,
	dreg_121,
	full_flag1,
	GND_port,
	clk_32_clk,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_34;
output 	q_b_33;
output 	q_b_35;
output 	q_b_32;
output 	q_b_28;
output 	q_b_24;
output 	q_b_29;
output 	q_b_25;
output 	q_b_30;
output 	q_b_26;
output 	q_b_31;
output 	q_b_27;
output 	q_b_20;
output 	q_b_16;
output 	q_b_21;
output 	q_b_17;
output 	q_b_22;
output 	q_b_18;
output 	q_b_23;
output 	q_b_19;
output 	q_b_12;
output 	q_b_8;
output 	q_b_13;
output 	q_b_9;
output 	q_b_14;
output 	q_b_10;
output 	q_b_15;
output 	q_b_11;
output 	q_b_4;
output 	q_b_0;
output 	q_b_5;
output 	q_b_1;
output 	q_b_6;
output 	q_b_2;
output 	q_b_7;
output 	q_b_3;
output 	septy_flag1;
output 	afull_flag1;
output 	aempty_flag1;
input 	dreg_1;
input 	dreg_11;
input 	dreg_12;
input 	dreg_13;
input 	dreg_14;
input 	dreg_15;
input 	dreg_16;
input 	dreg_17;
input 	dreg_18;
input 	dreg_19;
input 	dreg_110;
input 	altera_tse_reset_synchronizer_chain_out;
input 	altera_tse_reset_synchronizer_chain_out1;
output 	sav_flag1;
output 	empty_flag1;
input 	always5;
input 	dreg_111;
input 	dreg_112;
input 	dreg_113;
input 	dreg_114;
input 	dreg_115;
input 	dreg_116;
input 	dreg_117;
input 	dreg_118;
input 	dreg_119;
input 	dreg_120;
input 	dreg_121;
output 	full_flag1;
input 	GND_port;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_WRT|b_out[10]~q ;
wire \U_WRT|b_out[1]~q ;
wire \U_WRT|b_out[0]~q ;
wire \U_WRT|b_out[3]~q ;
wire \U_WRT|b_out[2]~q ;
wire \U_WRT|b_out[5]~q ;
wire \U_WRT|b_out[4]~q ;
wire \U_WRT|b_out[7]~q ;
wire \U_WRT|b_out[6]~q ;
wire \U_WRT|b_out[9]~q ;
wire \U_WRT|b_out[8]~q ;
wire \U_RD|b_out[10]~q ;
wire \U_RD|b_out[7]~q ;
wire \U_RD|b_out[6]~q ;
wire \U_RD|b_out[3]~q ;
wire \U_RD|b_out[2]~q ;
wire \U_RD|b_out[1]~q ;
wire \U_RD|b_out[0]~q ;
wire \U_RD|b_out[5]~q ;
wire \U_RD|b_out[4]~q ;
wire \U_RD|b_out[9]~q ;
wire \U_RD|b_out[8]~q ;
wire \U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[5].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ;
wire \U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ;
wire \U_RD|g_out[10]~q ;
wire \U_RD|g_out[9]~q ;
wire \U_RD|g_out[8]~q ;
wire \U_RD|g_out[7]~q ;
wire \U_RD|g_out[6]~q ;
wire \U_RD|g_out[5]~q ;
wire \U_RD|g_out[4]~q ;
wire \U_RD|g_out[3]~q ;
wire \U_RD|g_out[2]~q ;
wire \U_RD|g_out[1]~q ;
wire \U_RD|g_out[0]~q ;
wire \U_WRT|g_out[10]~q ;
wire \U_WRT|g_out[9]~q ;
wire \U_WRT|g_out[8]~q ;
wire \U_WRT|g_out[7]~q ;
wire \U_WRT|g_out[6]~q ;
wire \U_WRT|g_out[5]~q ;
wire \U_WRT|g_out[4]~q ;
wire \U_WRT|g_out[3]~q ;
wire \U_WRT|g_out[2]~q ;
wire \U_WRT|g_out[1]~q ;
wire \U_WRT|g_out[0]~q ;
wire \rd_b_wptr[10]~q ;
wire \ff_rd_binval[9]~7_combout ;
wire \rd_b_wptr[9]~q ;
wire \ff_rd_binval[8]~8_combout ;
wire \rd_b_wptr[8]~q ;
wire \ff_rd_binval[6]~5_combout ;
wire \rd_b_wptr[7]~q ;
wire \ff_rd_binval[6]~6_combout ;
wire \rd_b_wptr[6]~q ;
wire \ff_rd_binval[4]~0_combout ;
wire \rd_b_wptr[5]~q ;
wire \ff_rd_binval[4]~4_combout ;
wire \rd_b_wptr[4]~q ;
wire \ff_rd_binval[3]~2_combout ;
wire \rd_b_wptr[3]~q ;
wire \ff_rd_binval[1]~3_combout ;
wire \rd_b_wptr[2]~q ;
wire \ff_rd_binval[0]~1_combout ;
wire \rd_b_wptr[1]~q ;
wire \ff_rd_binval[0]~combout ;
wire \rd_b_wptr[0]~q ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~1_sumout ;
wire \ptr_wck_diff[10]~q ;
wire \LessThan2~0_combout ;
wire \Add0~5_sumout ;
wire \ptr_wck_diff[1]~q ;
wire \Add0~9_sumout ;
wire \ptr_wck_diff[0]~q ;
wire \LessThan2~1_combout ;
wire \Add0~13_sumout ;
wire \ptr_wck_diff[3]~q ;
wire \Add0~17_sumout ;
wire \ptr_wck_diff[2]~q ;
wire \LessThan2~2_combout ;
wire \LessThan2~3_combout ;
wire \Add0~21_sumout ;
wire \ptr_wck_diff[5]~q ;
wire \Add0~25_sumout ;
wire \ptr_wck_diff[4]~q ;
wire \LessThan2~4_combout ;
wire \LessThan2~5_combout ;
wire \Add0~29_sumout ;
wire \ptr_wck_diff[7]~q ;
wire \Add0~33_sumout ;
wire \ptr_wck_diff[6]~q ;
wire \LessThan2~6_combout ;
wire \LessThan2~7_combout ;
wire \LessThan2~8_combout ;
wire \Add0~37_sumout ;
wire \ptr_wck_diff[9]~q ;
wire \Add0~41_sumout ;
wire \ptr_wck_diff[8]~q ;
wire \septy_flag~0_combout ;
wire \septy_flag~1_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \septy_flag~2_combout ;
wire \septy_flag~3_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \LessThan0~3_combout ;
wire \LessThan0~4_combout ;
wire \LessThan0~5_combout ;
wire \LessThan0~6_combout ;
wire \LessThan0~7_combout ;
wire \LessThan0~8_combout ;
wire \afull_flag~0_combout ;
wire \afull_flag~1_combout ;
wire \afull_flag~2_combout ;
wire \afull_flag~3_combout ;
wire \afull_flag~4_combout ;
wire \afull_flag~5_combout ;
wire \wr_b_rptr[10]~q ;
wire \ff_wr_binval[9]~0_combout ;
wire \wr_b_rptr[9]~q ;
wire \ff_wr_binval[8]~1_combout ;
wire \wr_b_rptr[8]~q ;
wire \ff_wr_binval[6]~2_combout ;
wire \wr_b_rptr[7]~q ;
wire \ff_wr_binval[6]~3_combout ;
wire \wr_b_rptr[6]~q ;
wire \ff_wr_binval[4]~4_combout ;
wire \wr_b_rptr[5]~q ;
wire \ff_wr_binval[4]~8_combout ;
wire \wr_b_rptr[4]~q ;
wire \ff_wr_binval[3]~5_combout ;
wire \wr_b_rptr[3]~q ;
wire \ff_wr_binval[1]~6_combout ;
wire \wr_b_rptr[2]~q ;
wire \ff_wr_binval[0]~7_combout ;
wire \wr_b_rptr[1]~q ;
wire \ff_wr_binval[0]~combout ;
wire \wr_b_rptr[0]~q ;
wire \Add1~26 ;
wire \Add1~27 ;
wire \Add1~22 ;
wire \Add1~23 ;
wire \Add1~18 ;
wire \Add1~19 ;
wire \Add1~14 ;
wire \Add1~15 ;
wire \Add1~34 ;
wire \Add1~35 ;
wire \Add1~30 ;
wire \Add1~31 ;
wire \Add1~10 ;
wire \Add1~11 ;
wire \Add1~6 ;
wire \Add1~7 ;
wire \Add1~42 ;
wire \Add1~43 ;
wire \Add1~38 ;
wire \Add1~39 ;
wire \Add1~1_sumout ;
wire \ptr_rck_diff[10]~q ;
wire \Add1~5_sumout ;
wire \ptr_rck_diff[7]~q ;
wire \Add1~9_sumout ;
wire \ptr_rck_diff[6]~q ;
wire \Add1~13_sumout ;
wire \ptr_rck_diff[3]~q ;
wire \Add1~17_sumout ;
wire \ptr_rck_diff[2]~q ;
wire \Add1~21_sumout ;
wire \ptr_rck_diff[1]~q ;
wire \Add1~25_sumout ;
wire \ptr_rck_diff[0]~q ;
wire \LessThan3~0_combout ;
wire \Add1~29_sumout ;
wire \ptr_rck_diff[5]~q ;
wire \Add1~33_sumout ;
wire \ptr_rck_diff[4]~q ;
wire \LessThan3~1_combout ;
wire \LessThan3~2_combout ;
wire \LessThan3~3_combout ;
wire \LessThan3~4_combout ;
wire \Add1~37_sumout ;
wire \ptr_rck_diff[9]~q ;
wire \Add1~41_sumout ;
wire \ptr_rck_diff[8]~q ;
wire \aempty_flag~0_combout ;
wire \aempty_flag~1_combout ;
wire \aempty_flag~2_combout ;
wire \aempty_flag~3_combout ;
wire \aempty_flag~4_combout ;
wire \aempty_flag~5_combout ;
wire \LessThan4~0_combout ;
wire \LessThan4~1_combout ;
wire \LessThan4~2_combout ;
wire \LessThan4~3_combout ;
wire \LessThan4~4_combout ;
wire \sav_flag~0_combout ;
wire \sav_flag~1_combout ;
wire \Equal5~0_combout ;
wire \Equal5~1_combout ;
wire \Equal5~2_combout ;
wire \sav_flag~2_combout ;
wire \rden_reg~q ;
wire \empty_flag~0_combout ;
wire \empty_flag~1_combout ;
wire \empty_flag~2_combout ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;


IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_17 U_SYNC_4(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_16 U_SYNC_3(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out1),
	.dreg_1(\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_3|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.g_out_10(\U_WRT|g_out[10]~q ),
	.g_out_9(\U_WRT|g_out[9]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_15 U_SYNC_2(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_14 U_SYNC_1(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_11(\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_12(\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_13(\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_14(\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_15(\U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_16(\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_17(\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_18(\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_19(\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dreg_110(\U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.g_out_10(\U_RD|g_out[10]~q ),
	.g_out_9(\U_RD|g_out[9]~q ),
	.g_out_8(\U_RD|g_out[8]~q ),
	.g_out_7(\U_RD|g_out[7]~q ),
	.g_out_6(\U_RD|g_out[6]~q ),
	.g_out_5(\U_RD|g_out[5]~q ),
	.g_out_4(\U_RD|g_out[4]~q ),
	.g_out_3(\U_RD|g_out[3]~q ),
	.g_out_2(\U_RD|g_out[2]~q ),
	.g_out_1(\U_RD|g_out[1]~q ),
	.g_out_0(\U_RD|g_out[0]~q ),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_7 U_RD(
	.reset(altera_tse_reset_synchronizer_chain_out1),
	.b_out_10(\U_RD|b_out[10]~q ),
	.b_out_7(\U_RD|b_out[7]~q ),
	.b_out_6(\U_RD|b_out[6]~q ),
	.b_out_3(\U_RD|b_out[3]~q ),
	.b_out_2(\U_RD|b_out[2]~q ),
	.b_out_1(\U_RD|b_out[1]~q ),
	.b_out_0(\U_RD|b_out[0]~q ),
	.b_out_5(\U_RD|b_out[5]~q ),
	.b_out_4(\U_RD|b_out[4]~q ),
	.b_out_9(\U_RD|b_out[9]~q ),
	.b_out_8(\U_RD|b_out[8]~q ),
	.always5(always5),
	.g_out_10(\U_RD|g_out[10]~q ),
	.g_out_9(\U_RD|g_out[9]~q ),
	.g_out_8(\U_RD|g_out[8]~q ),
	.g_out_7(\U_RD|g_out[7]~q ),
	.g_out_6(\U_RD|g_out[6]~q ),
	.g_out_5(\U_RD|g_out[5]~q ),
	.g_out_4(\U_RD|g_out[4]~q ),
	.g_out_3(\U_RD|g_out[3]~q ),
	.g_out_2(\U_RD|g_out[2]~q ),
	.g_out_1(\U_RD|g_out[1]~q ),
	.g_out_0(\U_RD|g_out[0]~q ),
	.clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_tse_gray_cnt_8 U_WRT(
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.b_out_10(\U_WRT|b_out[10]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_9(\U_WRT|b_out[9]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.g_out_10(\U_WRT|g_out[10]~q ),
	.g_out_9(\U_WRT|g_out[9]~q ),
	.g_out_8(\U_WRT|g_out[8]~q ),
	.g_out_7(\U_WRT|g_out[7]~q ),
	.g_out_6(\U_WRT|g_out[6]~q ),
	.g_out_5(\U_WRT|g_out[5]~q ),
	.g_out_4(\U_WRT|g_out[4]~q ),
	.g_out_3(\U_WRT|g_out[3]~q ),
	.g_out_2(\U_WRT|g_out[2]~q ),
	.g_out_1(\U_WRT|g_out[1]~q ),
	.g_out_0(\U_WRT|g_out[0]~q ));

IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_3 U_RAM(
	.q_b_34(q_b_34),
	.q_b_33(q_b_33),
	.q_b_35(q_b_35),
	.q_b_32(q_b_32),
	.q_b_28(q_b_28),
	.q_b_24(q_b_24),
	.q_b_29(q_b_29),
	.q_b_25(q_b_25),
	.q_b_30(q_b_30),
	.q_b_26(q_b_26),
	.q_b_31(q_b_31),
	.q_b_27(q_b_27),
	.q_b_20(q_b_20),
	.q_b_16(q_b_16),
	.q_b_21(q_b_21),
	.q_b_17(q_b_17),
	.q_b_22(q_b_22),
	.q_b_18(q_b_18),
	.q_b_23(q_b_23),
	.q_b_19(q_b_19),
	.q_b_12(q_b_12),
	.q_b_8(q_b_8),
	.q_b_13(q_b_13),
	.q_b_9(q_b_9),
	.q_b_14(q_b_14),
	.q_b_10(q_b_10),
	.q_b_15(q_b_15),
	.q_b_11(q_b_11),
	.q_b_4(q_b_4),
	.q_b_0(q_b_0),
	.q_b_5(q_b_5),
	.q_b_1(q_b_1),
	.q_b_6(q_b_6),
	.q_b_2(q_b_2),
	.q_b_7(q_b_7),
	.q_b_3(q_b_3),
	.b_out_10(\U_WRT|b_out[10]~q ),
	.b_out_1(\U_WRT|b_out[1]~q ),
	.b_out_0(\U_WRT|b_out[0]~q ),
	.b_out_3(\U_WRT|b_out[3]~q ),
	.b_out_2(\U_WRT|b_out[2]~q ),
	.b_out_5(\U_WRT|b_out[5]~q ),
	.b_out_4(\U_WRT|b_out[4]~q ),
	.b_out_7(\U_WRT|b_out[7]~q ),
	.b_out_6(\U_WRT|b_out[6]~q ),
	.b_out_9(\U_WRT|b_out[9]~q ),
	.b_out_8(\U_WRT|b_out[8]~q ),
	.b_out_101(\U_RD|b_out[10]~q ),
	.b_out_71(\U_RD|b_out[7]~q ),
	.b_out_61(\U_RD|b_out[6]~q ),
	.b_out_31(\U_RD|b_out[3]~q ),
	.b_out_21(\U_RD|b_out[2]~q ),
	.b_out_11(\U_RD|b_out[1]~q ),
	.b_out_01(\U_RD|b_out[0]~q ),
	.b_out_51(\U_RD|b_out[5]~q ),
	.b_out_41(\U_RD|b_out[4]~q ),
	.b_out_91(\U_RD|b_out[9]~q ),
	.b_out_81(\U_RD|b_out[8]~q ),
	.GND_port(GND_port),
	.clk_32_clk(clk_32_clk),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

dffeas septy_flag(
	.clk(clk_32_clk),
	.d(\septy_flag~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(septy_flag1),
	.prn(vcc));
defparam septy_flag.is_wysiwyg = "true";
defparam septy_flag.power_up = "low";

dffeas afull_flag(
	.clk(clk_32_clk),
	.d(\afull_flag~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(afull_flag1),
	.prn(vcc));
defparam afull_flag.is_wysiwyg = "true";
defparam afull_flag.power_up = "low";

dffeas aempty_flag(
	.clk(mac_tx_clock_connection_clk),
	.d(\aempty_flag~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(aempty_flag1),
	.prn(vcc));
defparam aempty_flag.is_wysiwyg = "true";
defparam aempty_flag.power_up = "low";

dffeas sav_flag(
	.clk(mac_tx_clock_connection_clk),
	.d(\sav_flag~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sav_flag1),
	.prn(vcc));
defparam sav_flag.is_wysiwyg = "true";
defparam sav_flag.power_up = "low";

dffeas empty_flag(
	.clk(mac_tx_clock_connection_clk),
	.d(\empty_flag~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(empty_flag1),
	.prn(vcc));
defparam empty_flag.is_wysiwyg = "true";
defparam empty_flag.power_up = "low";

dffeas full_flag(
	.clk(clk_32_clk),
	.d(\LessThan1~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full_flag1),
	.prn(vcc));
defparam full_flag.is_wysiwyg = "true";
defparam full_flag.power_up = "low";

dffeas \rd_b_wptr[10] (
	.clk(clk_32_clk),
	.d(\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[10]~q ),
	.prn(vcc));
defparam \rd_b_wptr[10] .is_wysiwyg = "true";
defparam \rd_b_wptr[10] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[9]~7 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[9]~7 .extended_lut = "off";
defparam \ff_rd_binval[9]~7 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[9]~7 .shared_arith = "off";

dffeas \rd_b_wptr[9] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[9]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[9]~q ),
	.prn(vcc));
defparam \rd_b_wptr[9] .is_wysiwyg = "true";
defparam \rd_b_wptr[9] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[8]~8 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[8]~8 .extended_lut = "off";
defparam \ff_rd_binval[8]~8 .lut_mask = 64'h9696969696969696;
defparam \ff_rd_binval[8]~8 .shared_arith = "off";

dffeas \rd_b_wptr[8] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[8]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[8]~q ),
	.prn(vcc));
defparam \rd_b_wptr[8] .is_wysiwyg = "true";
defparam \rd_b_wptr[8] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[6]~5 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[6]~5 .extended_lut = "off";
defparam \ff_rd_binval[6]~5 .lut_mask = 64'h6996699669966996;
defparam \ff_rd_binval[6]~5 .shared_arith = "off";

dffeas \rd_b_wptr[7] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[6]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[7]~q ),
	.prn(vcc));
defparam \rd_b_wptr[7] .is_wysiwyg = "true";
defparam \rd_b_wptr[7] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[6]~6 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[6]~6 .extended_lut = "off";
defparam \ff_rd_binval[6]~6 .lut_mask = 64'h9669699696696996;
defparam \ff_rd_binval[6]~6 .shared_arith = "off";

dffeas \rd_b_wptr[6] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[6]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[6]~q ),
	.prn(vcc));
defparam \rd_b_wptr[6] .is_wysiwyg = "true";
defparam \rd_b_wptr[6] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[4]~0 (
	.dataa(!\U_SYNC_1|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_1|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_1|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[4]~0 .extended_lut = "off";
defparam \ff_rd_binval[4]~0 .lut_mask = 64'h6996966996696996;
defparam \ff_rd_binval[4]~0 .shared_arith = "off";

dffeas \rd_b_wptr[5] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[4]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[5]~q ),
	.prn(vcc));
defparam \rd_b_wptr[5] .is_wysiwyg = "true";
defparam \rd_b_wptr[5] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[4]~4 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[4]~4 .extended_lut = "off";
defparam \ff_rd_binval[4]~4 .lut_mask = 64'h6666666666666666;
defparam \ff_rd_binval[4]~4 .shared_arith = "off";

dffeas \rd_b_wptr[4] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[4]~q ),
	.prn(vcc));
defparam \rd_b_wptr[4] .is_wysiwyg = "true";
defparam \rd_b_wptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[3]~2 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[3]~2 .extended_lut = "off";
defparam \ff_rd_binval[3]~2 .lut_mask = 64'h9696969696969696;
defparam \ff_rd_binval[3]~2 .shared_arith = "off";

dffeas \rd_b_wptr[3] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[3]~q ),
	.prn(vcc));
defparam \rd_b_wptr[3] .is_wysiwyg = "true";
defparam \rd_b_wptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[1]~3 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[1]~3 .extended_lut = "off";
defparam \ff_rd_binval[1]~3 .lut_mask = 64'h6996699669966996;
defparam \ff_rd_binval[1]~3 .shared_arith = "off";

dffeas \rd_b_wptr[2] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[1]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[2]~q ),
	.prn(vcc));
defparam \rd_b_wptr[2] .is_wysiwyg = "true";
defparam \rd_b_wptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[0]~1 (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[0]~1 .extended_lut = "off";
defparam \ff_rd_binval[0]~1 .lut_mask = 64'h9669699696696996;
defparam \ff_rd_binval[0]~1 .shared_arith = "off";

dffeas \rd_b_wptr[1] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[0]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[1]~q ),
	.prn(vcc));
defparam \rd_b_wptr[1] .is_wysiwyg = "true";
defparam \rd_b_wptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_rd_binval[0] (
	.dataa(!\ff_rd_binval[4]~0_combout ),
	.datab(!\U_SYNC_1|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_1|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_1|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_1|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_1|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_rd_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_rd_binval[0] .extended_lut = "off";
defparam \ff_rd_binval[0] .lut_mask = 64'h6996966996696996;
defparam \ff_rd_binval[0] .shared_arith = "off";

dffeas \rd_b_wptr[0] (
	.clk(clk_32_clk),
	.d(\ff_rd_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_b_wptr[0]~q ),
	.prn(vcc));
defparam \rd_b_wptr[0] .is_wysiwyg = "true";
defparam \rd_b_wptr[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[0]~q ),
	.datad(!\U_WRT|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[1]~q ),
	.datad(!\U_WRT|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[2]~q ),
	.datad(!\U_WRT|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[3]~q ),
	.datad(!\U_WRT|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[4]~q ),
	.datad(!\U_WRT|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[5]~q ),
	.datad(!\U_WRT|b_out[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[6]~q ),
	.datad(!\U_WRT|b_out[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[7]~q ),
	.datad(!\U_WRT|b_out[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[8]~q ),
	.datad(!\U_WRT|b_out[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[9]~q ),
	.datad(!\U_WRT|b_out[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000F0FF00000FF0;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\rd_b_wptr[10]~q ),
	.datad(!\U_WRT|b_out[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000000000000FF0;
defparam \Add0~1 .shared_arith = "on";

dffeas \ptr_wck_diff[10] (
	.clk(clk_32_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[10]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[10] .is_wysiwyg = "true";
defparam \ptr_wck_diff[10] .power_up = "low";

cyclonev_lcell_comb \LessThan2~0 (
	.dataa(!dreg_1),
	.datab(!\ptr_wck_diff[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~0 .extended_lut = "off";
defparam \LessThan2~0 .lut_mask = 64'h6666666666666666;
defparam \LessThan2~0 .shared_arith = "off";

dffeas \ptr_wck_diff[1] (
	.clk(clk_32_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[1]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[1] .is_wysiwyg = "true";
defparam \ptr_wck_diff[1] .power_up = "low";

dffeas \ptr_wck_diff[0] (
	.clk(clk_32_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[0]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[0] .is_wysiwyg = "true";
defparam \ptr_wck_diff[0] .power_up = "low";

cyclonev_lcell_comb \LessThan2~1 (
	.dataa(!dreg_11),
	.datab(!dreg_12),
	.datac(!\ptr_wck_diff[1]~q ),
	.datad(!\ptr_wck_diff[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~1 .extended_lut = "off";
defparam \LessThan2~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan2~1 .shared_arith = "off";

dffeas \ptr_wck_diff[3] (
	.clk(clk_32_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[3]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[3] .is_wysiwyg = "true";
defparam \ptr_wck_diff[3] .power_up = "low";

dffeas \ptr_wck_diff[2] (
	.clk(clk_32_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[2]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[2] .is_wysiwyg = "true";
defparam \ptr_wck_diff[2] .power_up = "low";

cyclonev_lcell_comb \LessThan2~2 (
	.dataa(!dreg_13),
	.datab(!dreg_14),
	.datac(!\ptr_wck_diff[3]~q ),
	.datad(!\ptr_wck_diff[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~2 .extended_lut = "off";
defparam \LessThan2~2 .lut_mask = 64'h6996699669966996;
defparam \LessThan2~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~3 (
	.dataa(!dreg_13),
	.datab(!dreg_14),
	.datac(!\ptr_wck_diff[3]~q ),
	.datad(!\ptr_wck_diff[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~3 .extended_lut = "off";
defparam \LessThan2~3 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan2~3 .shared_arith = "off";

dffeas \ptr_wck_diff[5] (
	.clk(clk_32_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[5]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[5] .is_wysiwyg = "true";
defparam \ptr_wck_diff[5] .power_up = "low";

dffeas \ptr_wck_diff[4] (
	.clk(clk_32_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[4]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[4] .is_wysiwyg = "true";
defparam \ptr_wck_diff[4] .power_up = "low";

cyclonev_lcell_comb \LessThan2~4 (
	.dataa(!dreg_15),
	.datab(!dreg_16),
	.datac(!\ptr_wck_diff[5]~q ),
	.datad(!\ptr_wck_diff[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~4 .extended_lut = "off";
defparam \LessThan2~4 .lut_mask = 64'h6996699669966996;
defparam \LessThan2~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~5 (
	.dataa(!dreg_15),
	.datab(!dreg_16),
	.datac(!\ptr_wck_diff[5]~q ),
	.datad(!\ptr_wck_diff[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~5 .extended_lut = "off";
defparam \LessThan2~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan2~5 .shared_arith = "off";

dffeas \ptr_wck_diff[7] (
	.clk(clk_32_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[7]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[7] .is_wysiwyg = "true";
defparam \ptr_wck_diff[7] .power_up = "low";

dffeas \ptr_wck_diff[6] (
	.clk(clk_32_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[6]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[6] .is_wysiwyg = "true";
defparam \ptr_wck_diff[6] .power_up = "low";

cyclonev_lcell_comb \LessThan2~6 (
	.dataa(!dreg_17),
	.datab(!dreg_18),
	.datac(!\ptr_wck_diff[7]~q ),
	.datad(!\ptr_wck_diff[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~6 .extended_lut = "off";
defparam \LessThan2~6 .lut_mask = 64'h6996699669966996;
defparam \LessThan2~6 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~7 (
	.dataa(!\LessThan2~1_combout ),
	.datab(!\LessThan2~2_combout ),
	.datac(!\LessThan2~3_combout ),
	.datad(!\LessThan2~4_combout ),
	.datae(!\LessThan2~5_combout ),
	.dataf(!\LessThan2~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~7 .extended_lut = "off";
defparam \LessThan2~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \LessThan2~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~8 (
	.dataa(!dreg_17),
	.datab(!dreg_18),
	.datac(!\ptr_wck_diff[7]~q ),
	.datad(!\ptr_wck_diff[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~8 .extended_lut = "off";
defparam \LessThan2~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \LessThan2~8 .shared_arith = "off";

dffeas \ptr_wck_diff[9] (
	.clk(clk_32_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[9]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[9] .is_wysiwyg = "true";
defparam \ptr_wck_diff[9] .power_up = "low";

dffeas \ptr_wck_diff[8] (
	.clk(clk_32_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_wck_diff[8]~q ),
	.prn(vcc));
defparam \ptr_wck_diff[8] .is_wysiwyg = "true";
defparam \ptr_wck_diff[8] .power_up = "low";

cyclonev_lcell_comb \septy_flag~0 (
	.dataa(!dreg_19),
	.datab(!dreg_110),
	.datac(!\ptr_wck_diff[9]~q ),
	.datad(!\ptr_wck_diff[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\septy_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \septy_flag~0 .extended_lut = "off";
defparam \septy_flag~0 .lut_mask = 64'h6996699669966996;
defparam \septy_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \septy_flag~1 (
	.dataa(!dreg_19),
	.datab(!dreg_110),
	.datac(!\ptr_wck_diff[9]~q ),
	.datad(!\ptr_wck_diff[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\septy_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \septy_flag~1 .extended_lut = "off";
defparam \septy_flag~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \septy_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!dreg_11),
	.datab(!dreg_12),
	.datac(!dreg_13),
	.datad(!dreg_14),
	.datae(!dreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!dreg_17),
	.datab(!dreg_18),
	.datac(!dreg_19),
	.datad(!dreg_110),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \septy_flag~2 (
	.dataa(!dreg_16),
	.datab(!dreg_1),
	.datac(!\ptr_wck_diff[10]~q ),
	.datad(!\Equal1~0_combout ),
	.datae(!\Equal1~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\septy_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \septy_flag~2 .extended_lut = "off";
defparam \septy_flag~2 .lut_mask = 64'hB8FFFFFFB8FFFFFF;
defparam \septy_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \septy_flag~3 (
	.dataa(!\LessThan2~0_combout ),
	.datab(!\LessThan2~7_combout ),
	.datac(!\LessThan2~8_combout ),
	.datad(!\septy_flag~0_combout ),
	.datae(!\septy_flag~1_combout ),
	.dataf(!\septy_flag~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\septy_flag~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \septy_flag~3 .extended_lut = "off";
defparam \septy_flag~3 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \septy_flag~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\ptr_wck_diff[10]~q ),
	.datab(!\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h6666666666666666;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\ptr_wck_diff[1]~q ),
	.datab(!\ptr_wck_diff[0]~q ),
	.datac(!\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!\ptr_wck_diff[3]~q ),
	.datab(!\ptr_wck_diff[2]~q ),
	.datac(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h6996699669966996;
defparam \LessThan0~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~3 (
	.dataa(!\ptr_wck_diff[3]~q ),
	.datab(!\ptr_wck_diff[2]~q ),
	.datac(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~3 .extended_lut = "off";
defparam \LessThan0~3 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~4 (
	.dataa(!\ptr_wck_diff[5]~q ),
	.datab(!\ptr_wck_diff[4]~q ),
	.datac(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~4 .extended_lut = "off";
defparam \LessThan0~4 .lut_mask = 64'h6996699669966996;
defparam \LessThan0~4 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~5 (
	.dataa(!\ptr_wck_diff[5]~q ),
	.datab(!\ptr_wck_diff[4]~q ),
	.datac(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~5 .extended_lut = "off";
defparam \LessThan0~5 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~6 (
	.dataa(!\ptr_wck_diff[7]~q ),
	.datab(!\ptr_wck_diff[6]~q ),
	.datac(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~6 .extended_lut = "off";
defparam \LessThan0~6 .lut_mask = 64'h6996699669966996;
defparam \LessThan0~6 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~7 (
	.dataa(!\LessThan0~1_combout ),
	.datab(!\LessThan0~2_combout ),
	.datac(!\LessThan0~3_combout ),
	.datad(!\LessThan0~4_combout ),
	.datae(!\LessThan0~5_combout ),
	.dataf(!\LessThan0~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~7 .extended_lut = "off";
defparam \LessThan0~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \LessThan0~7 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~8 (
	.dataa(!\ptr_wck_diff[7]~q ),
	.datab(!\ptr_wck_diff[6]~q ),
	.datac(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~8 .extended_lut = "off";
defparam \LessThan0~8 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~8 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~0 (
	.dataa(!\ptr_wck_diff[9]~q ),
	.datab(!\ptr_wck_diff[8]~q ),
	.datac(!\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~0 .extended_lut = "off";
defparam \afull_flag~0 .lut_mask = 64'h6996699669966996;
defparam \afull_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~1 (
	.dataa(!\ptr_wck_diff[9]~q ),
	.datab(!\ptr_wck_diff[8]~q ),
	.datac(!\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~1 .extended_lut = "off";
defparam \afull_flag~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \afull_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~2 (
	.dataa(!\U_SYNC_2|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_2|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~2 .extended_lut = "off";
defparam \afull_flag~2 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \afull_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~3 (
	.dataa(!\U_SYNC_2|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_2|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_2|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~3 .extended_lut = "off";
defparam \afull_flag~3 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \afull_flag~3 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~4 (
	.dataa(!\ptr_wck_diff[10]~q ),
	.datab(!\U_SYNC_2|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_2|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\afull_flag~2_combout ),
	.datae(!\afull_flag~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~4 .extended_lut = "off";
defparam \afull_flag~4 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \afull_flag~4 .shared_arith = "off";

cyclonev_lcell_comb \afull_flag~5 (
	.dataa(!\LessThan0~0_combout ),
	.datab(!\LessThan0~7_combout ),
	.datac(!\LessThan0~8_combout ),
	.datad(!\afull_flag~0_combout ),
	.datae(!\afull_flag~1_combout ),
	.dataf(!\afull_flag~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\afull_flag~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \afull_flag~5 .extended_lut = "off";
defparam \afull_flag~5 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \afull_flag~5 .shared_arith = "off";

dffeas \wr_b_rptr[10] (
	.clk(mac_tx_clock_connection_clk),
	.d(\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[10]~q ),
	.prn(vcc));
defparam \wr_b_rptr[10] .is_wysiwyg = "true";
defparam \wr_b_rptr[10] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[9]~0 (
	.dataa(!\U_SYNC_3|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_3|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[9]~0 .extended_lut = "off";
defparam \ff_wr_binval[9]~0 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[9]~0 .shared_arith = "off";

dffeas \wr_b_rptr[9] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[9]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[9]~q ),
	.prn(vcc));
defparam \wr_b_rptr[9] .is_wysiwyg = "true";
defparam \wr_b_rptr[9] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[8]~1 (
	.dataa(!\ff_wr_binval[9]~0_combout ),
	.datab(!\U_SYNC_3|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[8]~1 .extended_lut = "off";
defparam \ff_wr_binval[8]~1 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[8]~1 .shared_arith = "off";

dffeas \wr_b_rptr[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[8]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[8]~q ),
	.prn(vcc));
defparam \wr_b_rptr[8] .is_wysiwyg = "true";
defparam \wr_b_rptr[8] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[6]~2 (
	.dataa(!\ff_wr_binval[8]~1_combout ),
	.datab(!\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[6]~2 .extended_lut = "off";
defparam \ff_wr_binval[6]~2 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[6]~2 .shared_arith = "off";

dffeas \wr_b_rptr[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[6]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[7]~q ),
	.prn(vcc));
defparam \wr_b_rptr[7] .is_wysiwyg = "true";
defparam \wr_b_rptr[7] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[6]~3 (
	.dataa(!\ff_wr_binval[6]~2_combout ),
	.datab(!\U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[6]~3 .extended_lut = "off";
defparam \ff_wr_binval[6]~3 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[6]~3 .shared_arith = "off";

dffeas \wr_b_rptr[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[6]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[6]~q ),
	.prn(vcc));
defparam \wr_b_rptr[6] .is_wysiwyg = "true";
defparam \wr_b_rptr[6] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[4]~4 (
	.dataa(!\ff_wr_binval[8]~1_combout ),
	.datab(!\U_SYNC_3|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[4]~4 .extended_lut = "off";
defparam \ff_wr_binval[4]~4 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[4]~4 .shared_arith = "off";

dffeas \wr_b_rptr[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[4]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[5]~q ),
	.prn(vcc));
defparam \wr_b_rptr[5] .is_wysiwyg = "true";
defparam \wr_b_rptr[5] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[4]~8 (
	.dataa(!\ff_wr_binval[4]~4_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[4]~8 .extended_lut = "off";
defparam \ff_wr_binval[4]~8 .lut_mask = 64'h6666666666666666;
defparam \ff_wr_binval[4]~8 .shared_arith = "off";

dffeas \wr_b_rptr[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[4]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[4]~q ),
	.prn(vcc));
defparam \wr_b_rptr[4] .is_wysiwyg = "true";
defparam \wr_b_rptr[4] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[3]~5 (
	.dataa(!\ff_wr_binval[4]~4_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[3]~5 .extended_lut = "off";
defparam \ff_wr_binval[3]~5 .lut_mask = 64'h9696969696969696;
defparam \ff_wr_binval[3]~5 .shared_arith = "off";

dffeas \wr_b_rptr[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[3]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[3]~q ),
	.prn(vcc));
defparam \wr_b_rptr[3] .is_wysiwyg = "true";
defparam \wr_b_rptr[3] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[1]~6 (
	.dataa(!\ff_wr_binval[4]~4_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[1]~6 .extended_lut = "off";
defparam \ff_wr_binval[1]~6 .lut_mask = 64'h6996699669966996;
defparam \ff_wr_binval[1]~6 .shared_arith = "off";

dffeas \wr_b_rptr[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[1]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[2]~q ),
	.prn(vcc));
defparam \wr_b_rptr[2] .is_wysiwyg = "true";
defparam \wr_b_rptr[2] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0]~7 (
	.dataa(!\ff_wr_binval[4]~4_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0]~7 .extended_lut = "off";
defparam \ff_wr_binval[0]~7 .lut_mask = 64'h9669699696696996;
defparam \ff_wr_binval[0]~7 .shared_arith = "off";

dffeas \wr_b_rptr[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[0]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[1]~q ),
	.prn(vcc));
defparam \wr_b_rptr[1] .is_wysiwyg = "true";
defparam \wr_b_rptr[1] .power_up = "low";

cyclonev_lcell_comb \ff_wr_binval[0] (
	.dataa(!\ff_wr_binval[4]~4_combout ),
	.datab(!\U_SYNC_3|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_3|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_3|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\U_SYNC_3|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.dataf(!\U_SYNC_3|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ff_wr_binval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ff_wr_binval[0] .extended_lut = "off";
defparam \ff_wr_binval[0] .lut_mask = 64'h6996966996696996;
defparam \ff_wr_binval[0] .shared_arith = "off";

dffeas \wr_b_rptr[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\ff_wr_binval[0]~combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wr_b_rptr[0]~q ),
	.prn(vcc));
defparam \wr_b_rptr[0] .is_wysiwyg = "true";
defparam \wr_b_rptr[0] .power_up = "low";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[0]~q ),
	.datad(!\U_RD|b_out[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout(\Add1~27 ));
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~25 .shared_arith = "on";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[1]~q ),
	.datad(!\U_RD|b_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(\Add1~27 ),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout(\Add1~23 ));
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~21 .shared_arith = "on";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[2]~q ),
	.datad(!\U_RD|b_out[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(\Add1~23 ),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout(\Add1~19 ));
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~17 .shared_arith = "on";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[3]~q ),
	.datad(!\U_RD|b_out[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(\Add1~19 ),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout(\Add1~15 ));
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~13 .shared_arith = "on";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[4]~q ),
	.datad(!\U_RD|b_out[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(\Add1~15 ),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout(\Add1~35 ));
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~33 .shared_arith = "on";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[5]~q ),
	.datad(!\U_RD|b_out[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(\Add1~35 ),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout(\Add1~31 ));
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~29 .shared_arith = "on";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[6]~q ),
	.datad(!\U_RD|b_out[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(\Add1~31 ),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout(\Add1~11 ));
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~9 .shared_arith = "on";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[7]~q ),
	.datad(!\U_RD|b_out[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(\Add1~11 ),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout(\Add1~7 ));
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~5 .shared_arith = "on";

cyclonev_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[8]~q ),
	.datad(!\U_RD|b_out[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(\Add1~7 ),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout(\Add1~43 ));
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~41 .shared_arith = "on";

cyclonev_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[9]~q ),
	.datad(!\U_RD|b_out[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(\Add1~43 ),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout(\Add1~39 ));
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add1~37 .shared_arith = "on";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\wr_b_rptr[10]~q ),
	.datad(!\U_RD|b_out[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(\Add1~39 ),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000000000000FF0;
defparam \Add1~1 .shared_arith = "on";

dffeas \ptr_rck_diff[10] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[10]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[10] .is_wysiwyg = "true";
defparam \ptr_rck_diff[10] .power_up = "low";

dffeas \ptr_rck_diff[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[7]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[7] .is_wysiwyg = "true";
defparam \ptr_rck_diff[7] .power_up = "low";

dffeas \ptr_rck_diff[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[6]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[6] .is_wysiwyg = "true";
defparam \ptr_rck_diff[6] .power_up = "low";

dffeas \ptr_rck_diff[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[3]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[3] .is_wysiwyg = "true";
defparam \ptr_rck_diff[3] .power_up = "low";

dffeas \ptr_rck_diff[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[2]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[2] .is_wysiwyg = "true";
defparam \ptr_rck_diff[2] .power_up = "low";

dffeas \ptr_rck_diff[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[1]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[1] .is_wysiwyg = "true";
defparam \ptr_rck_diff[1] .power_up = "low";

dffeas \ptr_rck_diff[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[0]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[0] .is_wysiwyg = "true";
defparam \ptr_rck_diff[0] .power_up = "low";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!\ptr_rck_diff[1]~q ),
	.datab(!\U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[0]~q ),
	.datad(!\U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \LessThan3~0 .shared_arith = "off";

dffeas \ptr_rck_diff[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[5]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[5] .is_wysiwyg = "true";
defparam \ptr_rck_diff[5] .power_up = "low";

dffeas \ptr_rck_diff[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[4]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[4] .is_wysiwyg = "true";
defparam \ptr_rck_diff[4] .power_up = "low";

cyclonev_lcell_comb \LessThan3~1 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[4]~q ),
	.datad(!\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~1 .extended_lut = "off";
defparam \LessThan3~1 .lut_mask = 64'h6996699669966996;
defparam \LessThan3~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~2 (
	.dataa(!\ptr_rck_diff[3]~q ),
	.datab(!\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[2]~q ),
	.datad(!\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\LessThan3~0_combout ),
	.dataf(!\LessThan3~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~2 .extended_lut = "off";
defparam \LessThan3~2 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \LessThan3~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~3 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[4]~q ),
	.datad(!\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~3 .extended_lut = "off";
defparam \LessThan3~3 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \LessThan3~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~4 (
	.dataa(!\ptr_rck_diff[7]~q ),
	.datab(!\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[6]~q ),
	.datad(!\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(!\LessThan3~2_combout ),
	.dataf(!\LessThan3~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~4 .extended_lut = "off";
defparam \LessThan3~4 .lut_mask = 64'hFFFFFFFFFFFFFBFF;
defparam \LessThan3~4 .shared_arith = "off";

dffeas \ptr_rck_diff[9] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~37_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[9]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[9] .is_wysiwyg = "true";
defparam \ptr_rck_diff[9] .power_up = "low";

dffeas \ptr_rck_diff[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add1~41_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ptr_rck_diff[8]~q ),
	.prn(vcc));
defparam \ptr_rck_diff[8] .is_wysiwyg = "true";
defparam \ptr_rck_diff[8] .power_up = "low";

cyclonev_lcell_comb \aempty_flag~0 (
	.dataa(!\ptr_rck_diff[9]~q ),
	.datab(!\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[8]~q ),
	.datad(!\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~0 .extended_lut = "off";
defparam \aempty_flag~0 .lut_mask = 64'h6996699669966996;
defparam \aempty_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~1 (
	.dataa(!\ptr_rck_diff[9]~q ),
	.datab(!\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\ptr_rck_diff[8]~q ),
	.datad(!\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~1 .extended_lut = "off";
defparam \aempty_flag~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \aempty_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~2 (
	.dataa(!\U_SYNC_4|sync[3].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_4|sync[2].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_4|sync[1].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[0].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~2 .extended_lut = "off";
defparam \aempty_flag~2 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \aempty_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~3 (
	.dataa(!\U_SYNC_4|sync[9].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_4|sync[8].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\U_SYNC_4|sync[7].u|std_sync_no_cut|dreg[1]~q ),
	.datad(!\U_SYNC_4|sync[6].u|std_sync_no_cut|dreg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~3 .extended_lut = "off";
defparam \aempty_flag~3 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \aempty_flag~3 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~4 (
	.dataa(!\U_SYNC_4|sync[5].u|std_sync_no_cut|dreg[1]~q ),
	.datab(!\U_SYNC_4|sync[4].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\aempty_flag~2_combout ),
	.datad(!\aempty_flag~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~4 .extended_lut = "off";
defparam \aempty_flag~4 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \aempty_flag~4 .shared_arith = "off";

cyclonev_lcell_comb \aempty_flag~5 (
	.dataa(!\ptr_rck_diff[10]~q ),
	.datab(!\U_SYNC_4|sync[10].u|std_sync_no_cut|dreg[1]~q ),
	.datac(!\LessThan3~4_combout ),
	.datad(!\aempty_flag~0_combout ),
	.datae(!\aempty_flag~1_combout ),
	.dataf(!\aempty_flag~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\aempty_flag~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \aempty_flag~5 .extended_lut = "off";
defparam \aempty_flag~5 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \aempty_flag~5 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~0 (
	.dataa(!\ptr_rck_diff[1]~q ),
	.datab(!\ptr_rck_diff[0]~q ),
	.datac(!dreg_116),
	.datad(!dreg_117),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~0 .extended_lut = "off";
defparam \LessThan4~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \LessThan4~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~1 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\ptr_rck_diff[4]~q ),
	.datac(!dreg_118),
	.datad(!dreg_119),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~1 .extended_lut = "off";
defparam \LessThan4~1 .lut_mask = 64'h6996699669966996;
defparam \LessThan4~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~2 (
	.dataa(!\ptr_rck_diff[3]~q ),
	.datab(!\ptr_rck_diff[2]~q ),
	.datac(!dreg_114),
	.datad(!dreg_115),
	.datae(!\LessThan4~0_combout ),
	.dataf(!\LessThan4~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~2 .extended_lut = "off";
defparam \LessThan4~2 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \LessThan4~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~3 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\ptr_rck_diff[4]~q ),
	.datac(!dreg_118),
	.datad(!dreg_119),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~3 .extended_lut = "off";
defparam \LessThan4~3 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \LessThan4~3 .shared_arith = "off";

cyclonev_lcell_comb \LessThan4~4 (
	.dataa(!\ptr_rck_diff[7]~q ),
	.datab(!\ptr_rck_diff[6]~q ),
	.datac(!dreg_112),
	.datad(!dreg_113),
	.datae(!\LessThan4~2_combout ),
	.dataf(!\LessThan4~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan4~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan4~4 .extended_lut = "off";
defparam \LessThan4~4 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \LessThan4~4 .shared_arith = "off";

cyclonev_lcell_comb \sav_flag~0 (
	.dataa(!\ptr_rck_diff[9]~q ),
	.datab(!\ptr_rck_diff[8]~q ),
	.datac(!dreg_120),
	.datad(!dreg_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~0 .extended_lut = "off";
defparam \sav_flag~0 .lut_mask = 64'h6996699669966996;
defparam \sav_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \sav_flag~1 (
	.dataa(!\ptr_rck_diff[9]~q ),
	.datab(!\ptr_rck_diff[8]~q ),
	.datac(!dreg_120),
	.datad(!dreg_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~1 .extended_lut = "off";
defparam \sav_flag~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \sav_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~0 (
	.dataa(!dreg_116),
	.datab(!dreg_117),
	.datac(!dreg_114),
	.datad(!dreg_115),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~0 .extended_lut = "off";
defparam \Equal5~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~1 (
	.dataa(!dreg_112),
	.datab(!dreg_113),
	.datac(!dreg_120),
	.datad(!dreg_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~1 .extended_lut = "off";
defparam \Equal5~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal5~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal5~2 (
	.dataa(!dreg_118),
	.datab(!dreg_119),
	.datac(!dreg_111),
	.datad(!\Equal5~0_combout ),
	.datae(!\Equal5~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal5~2 .extended_lut = "off";
defparam \Equal5~2 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \Equal5~2 .shared_arith = "off";

cyclonev_lcell_comb \sav_flag~2 (
	.dataa(!\ptr_rck_diff[10]~q ),
	.datab(!dreg_111),
	.datac(!\LessThan4~4_combout ),
	.datad(!\sav_flag~0_combout ),
	.datae(!\sav_flag~1_combout ),
	.dataf(!\Equal5~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sav_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sav_flag~2 .extended_lut = "off";
defparam \sav_flag~2 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \sav_flag~2 .shared_arith = "off";

dffeas rden_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(always5),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rden_reg~q ),
	.prn(vcc));
defparam rden_reg.is_wysiwyg = "true";
defparam rden_reg.power_up = "low";

cyclonev_lcell_comb \empty_flag~0 (
	.dataa(!\ptr_rck_diff[10]~q ),
	.datab(!\ptr_rck_diff[9]~q ),
	.datac(!\ptr_rck_diff[8]~q ),
	.datad(!\ptr_rck_diff[7]~q ),
	.datae(!\ptr_rck_diff[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~0 .extended_lut = "off";
defparam \empty_flag~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \empty_flag~0 .shared_arith = "off";

cyclonev_lcell_comb \empty_flag~1 (
	.dataa(!\ptr_rck_diff[4]~q ),
	.datab(!\ptr_rck_diff[3]~q ),
	.datac(!\ptr_rck_diff[2]~q ),
	.datad(!\ptr_rck_diff[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~1 .extended_lut = "off";
defparam \empty_flag~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \empty_flag~1 .shared_arith = "off";

cyclonev_lcell_comb \empty_flag~2 (
	.dataa(!\ptr_rck_diff[5]~q ),
	.datab(!\ptr_rck_diff[0]~q ),
	.datac(!\rden_reg~q ),
	.datad(!\empty_flag~0_combout ),
	.datae(!\empty_flag~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\empty_flag~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \empty_flag~2 .extended_lut = "off";
defparam \empty_flag~2 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \empty_flag~2 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!\ptr_wck_diff[10]~q ),
	.datab(!\ptr_wck_diff[9]~q ),
	.datac(!\ptr_wck_diff[8]~q ),
	.datad(!\ptr_wck_diff[7]~q ),
	.datae(!\ptr_wck_diff[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\ptr_wck_diff[5]~q ),
	.datab(!\ptr_wck_diff[4]~q ),
	.datac(!\ptr_wck_diff[3]~q ),
	.datad(!\ptr_wck_diff[2]~q ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan1~1 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_14 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	g_out_10;
input 	g_out_9;
input 	g_out_8;
input 	g_out_7;
input 	g_out_6;
input 	g_out_5;
input 	g_out_4;
input 	g_out_3;
input 	g_out_2;
input 	g_out_1;
input 	g_out_0;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_184 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.g_out_10(g_out_10),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_193 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.g_out_9(g_out_9),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_192 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.g_out_8(g_out_8),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_191 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.g_out_7(g_out_7),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_190 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.g_out_6(g_out_6),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_189 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.g_out_5(g_out_5),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_188 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.g_out_4(g_out_4),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_187 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.g_out_3(g_out_3),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_186 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.g_out_2(g_out_2),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_185 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.g_out_1(g_out_1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_183 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.g_out_0(g_out_0),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_183 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_0,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_0;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_183 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_0),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_183 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_184 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_10,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_10;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_184 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_10),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_184 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_185 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_185 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_185 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_186 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_2,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_2;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_186 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_2),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_186 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_187 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_3,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_3;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_187 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_3),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_187 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_188 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_4,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_4;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_188 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_4),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_188 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_189 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_5,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_5;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_189 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_5),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_189 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_190 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_6,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_6;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_190 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_6),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_190 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_191 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_7,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_7;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_191 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_7),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_191 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_192 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_8,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_8;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_192 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_8),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_192 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_193 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_9,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_9;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_193 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_9),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_193 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_15 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_195 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_204 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_203 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_202 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_201 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_200 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_199 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_198 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_197 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_196 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.clk_32_clk(clk_32_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_194 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.clk_32_clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_194 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_194 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_194 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_195 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_195 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_195 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_196 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_196 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_196 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_197 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_197 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_197 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_198 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_198 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_198 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_199 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_199 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_199 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_200 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_200 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_200 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_201 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_201 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_201 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_202 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_202 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_202 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_203 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_203 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_203 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_204 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	clk_32_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	clk_32_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_204 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(clk_32_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_204 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_16 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	g_out_10;
input 	g_out_9;
input 	g_out_8;
input 	g_out_7;
input 	g_out_6;
input 	g_out_5;
input 	g_out_4;
input 	g_out_3;
input 	g_out_2;
input 	g_out_1;
input 	g_out_0;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_206 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.g_out_10(g_out_10),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_215 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.g_out_9(g_out_9),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_214 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.g_out_8(g_out_8),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_213 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.g_out_7(g_out_7),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_212 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.g_out_6(g_out_6),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_211 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.g_out_5(g_out_5),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_210 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.g_out_4(g_out_4),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_209 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.g_out_3(g_out_3),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_208 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.g_out_2(g_out_2),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_207 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.g_out_1(g_out_1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_205 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.g_out_0(g_out_0),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_205 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_0,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_0;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_205 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_0),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_205 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_206 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_10,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_10;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_206 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_10),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_206 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_207 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_207 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_207 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_208 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_2,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_2;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_208 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_2),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_208 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_209 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_3,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_3;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_209 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_3),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_209 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_210 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_4,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_4;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_210 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_4),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_210 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_211 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_5,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_5;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_211 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_5),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_211 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_212 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_6,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_6;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_212 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_6),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_212 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_213 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_7,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_7;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_213 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_7),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_213 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_214 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_8,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_8;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_214 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_8),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_214 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_215 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	g_out_9,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	g_out_9;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_215 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.din(g_out_9),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_215 (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_bundle_17 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	dreg_11,
	dreg_12,
	dreg_13,
	dreg_14,
	dreg_15,
	dreg_16,
	dreg_17,
	dreg_18,
	dreg_19,
	dreg_110,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
output 	dreg_11;
output 	dreg_12;
output 	dreg_13;
output 	dreg_14;
output 	dreg_15;
output 	dreg_16;
output 	dreg_17;
output 	dreg_18;
output 	dreg_19;
output 	dreg_110;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_217 \sync[10].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_226 \sync[9].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_19),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_225 \sync[8].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_110),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_224 \sync[7].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_11),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_223 \sync[6].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_12),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_222 \sync[5].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_17),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_221 \sync[4].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_18),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_220 \sync[3].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_13),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_219 \sync[2].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_14),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_218 \sync[1].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_15),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_216 \sync[0].u (
	.altera_tse_reset_synchronizer_chain_out(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_16),
	.mac_tx_clock_connection_clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_216 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_216 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_216 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_217 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_217 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_217 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_218 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_218 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_218 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_219 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_219 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_219 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_220 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_220 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_220 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_221 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_221 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_221 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_222 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_222 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_222 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_223 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_223 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_223 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_224 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_224 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_224 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_225 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_225 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_225 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_eth_tse_std_synchronizer_226 (
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	dreg_1;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altera_std_synchronizer_nocut_226 std_sync_no_cut(
	.reset_n(altera_tse_reset_synchronizer_chain_out),
	.dreg_1(dreg_1),
	.clk(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altera_std_synchronizer_nocut_226 (
	reset_n,
	dreg_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~0_combout ;
wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

cyclonev_lcell_comb \din_s1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\din_s1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \din_s1~0 .extended_lut = "off";
defparam \din_s1~0 .lut_mask = 64'h0000000000000000;
defparam \din_s1~0 .shared_arith = "off";

dffeas din_s1(
	.clk(clk),
	.d(\din_s1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_3 (
	q_b_34,
	q_b_33,
	q_b_35,
	q_b_32,
	q_b_28,
	q_b_24,
	q_b_29,
	q_b_25,
	q_b_30,
	q_b_26,
	q_b_31,
	q_b_27,
	q_b_20,
	q_b_16,
	q_b_21,
	q_b_17,
	q_b_22,
	q_b_18,
	q_b_23,
	q_b_19,
	q_b_12,
	q_b_8,
	q_b_13,
	q_b_9,
	q_b_14,
	q_b_10,
	q_b_15,
	q_b_11,
	q_b_4,
	q_b_0,
	q_b_5,
	q_b_1,
	q_b_6,
	q_b_2,
	q_b_7,
	q_b_3,
	b_out_10,
	b_out_1,
	b_out_0,
	b_out_3,
	b_out_2,
	b_out_5,
	b_out_4,
	b_out_7,
	b_out_6,
	b_out_9,
	b_out_8,
	b_out_101,
	b_out_71,
	b_out_61,
	b_out_31,
	b_out_21,
	b_out_11,
	b_out_01,
	b_out_51,
	b_out_41,
	b_out_91,
	b_out_81,
	GND_port,
	clk_32_clk,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_34;
output 	q_b_33;
output 	q_b_35;
output 	q_b_32;
output 	q_b_28;
output 	q_b_24;
output 	q_b_29;
output 	q_b_25;
output 	q_b_30;
output 	q_b_26;
output 	q_b_31;
output 	q_b_27;
output 	q_b_20;
output 	q_b_16;
output 	q_b_21;
output 	q_b_17;
output 	q_b_22;
output 	q_b_18;
output 	q_b_23;
output 	q_b_19;
output 	q_b_12;
output 	q_b_8;
output 	q_b_13;
output 	q_b_9;
output 	q_b_14;
output 	q_b_10;
output 	q_b_15;
output 	q_b_11;
output 	q_b_4;
output 	q_b_0;
output 	q_b_5;
output 	q_b_1;
output 	q_b_6;
output 	q_b_2;
output 	q_b_7;
output 	q_b_3;
input 	b_out_10;
input 	b_out_1;
input 	b_out_0;
input 	b_out_3;
input 	b_out_2;
input 	b_out_5;
input 	b_out_4;
input 	b_out_7;
input 	b_out_6;
input 	b_out_9;
input 	b_out_8;
input 	b_out_101;
input 	b_out_71;
input 	b_out_61;
input 	b_out_31;
input 	b_out_21;
input 	b_out_11;
input 	b_out_01;
input 	b_out_51;
input 	b_out_41;
input 	b_out_91;
input 	b_out_81;
input 	GND_port;
input 	clk_32_clk;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_5 altsyncram_component(
	.q_b({q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_35,q_b_34,q_b_33,q_b_32,q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,
q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({b_out_10,b_out_9,b_out_8,b_out_7,b_out_6,b_out_5,b_out_4,b_out_3,b_out_2,b_out_1,b_out_0}),
	.address_b({b_out_101,b_out_91,b_out_81,b_out_71,b_out_61,b_out_51,b_out_41,b_out_31,b_out_21,b_out_11,b_out_01}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,GND_port,gnd,gnd,gnd}),
	.clock0(clk_32_clk),
	.clock1(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altsyncram_5 (
	q_b,
	address_a,
	address_b,
	data_a,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	[10:0] address_a;
input 	[10:0] address_b;
input 	[39:0] data_a;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_3ao1 auto_generated(
	.q_b({q_b[35],q_b[34],q_b[33],q_b[32],q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.data_a({data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3],data_a[3]}),
	.clock0(clock0),
	.clock1(clock1));

endmodule

module IoTOctopus_QSYS_altsyncram_3ao1 (
	q_b,
	address_a,
	address_b,
	data_a,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[35:0] q_b;
input 	[10:0] address_a;
input 	[10:0] address_b;
input 	[35:0] data_a;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[34] = ram_block1a34_PORTBDATAOUT_bus[0];

assign q_b[33] = ram_block1a33_PORTBDATAOUT_bus[0];

assign q_b[35] = ram_block1a35_PORTBDATAOUT_bus[0];

assign q_b[32] = ram_block1a32_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a34(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 11;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 2047;
defparam ram_block1a34.port_a_logical_ram_depth = 2048;
defparam ram_block1a34.port_a_logical_ram_width = 36;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 11;
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "none";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 2047;
defparam ram_block1a34.port_b_logical_ram_depth = 2048;
defparam ram_block1a34.port_b_logical_ram_width = 36;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";

cyclonev_ram_block ram_block1a33(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 11;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 2047;
defparam ram_block1a33.port_a_logical_ram_depth = 2048;
defparam ram_block1a33.port_a_logical_ram_width = 36;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 11;
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "none";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 2047;
defparam ram_block1a33.port_b_logical_ram_depth = 2048;
defparam ram_block1a33.port_b_logical_ram_width = 36;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";

cyclonev_ram_block ram_block1a35(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 11;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 2047;
defparam ram_block1a35.port_a_logical_ram_depth = 2048;
defparam ram_block1a35.port_a_logical_ram_width = 36;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 11;
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "none";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 2047;
defparam ram_block1a35.port_b_logical_ram_depth = 2048;
defparam ram_block1a35.port_b_logical_ram_width = 36;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";

cyclonev_ram_block ram_block1a32(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 11;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 2047;
defparam ram_block1a32.port_a_logical_ram_depth = 2048;
defparam ram_block1a32.port_a_logical_ram_width = 36;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 11;
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "none";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 2047;
defparam ram_block1a32.port_b_logical_ram_depth = 2048;
defparam ram_block1a32.port_b_logical_ram_width = 36;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 11;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 2047;
defparam ram_block1a28.port_a_logical_ram_depth = 2048;
defparam ram_block1a28.port_a_logical_ram_width = 36;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 11;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 2047;
defparam ram_block1a28.port_b_logical_ram_depth = 2048;
defparam ram_block1a28.port_b_logical_ram_width = 36;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 11;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 2047;
defparam ram_block1a24.port_a_logical_ram_depth = 2048;
defparam ram_block1a24.port_a_logical_ram_width = 36;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 11;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 2047;
defparam ram_block1a24.port_b_logical_ram_depth = 2048;
defparam ram_block1a24.port_b_logical_ram_width = 36;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 11;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 2047;
defparam ram_block1a29.port_a_logical_ram_depth = 2048;
defparam ram_block1a29.port_a_logical_ram_width = 36;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 11;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 2047;
defparam ram_block1a29.port_b_logical_ram_depth = 2048;
defparam ram_block1a29.port_b_logical_ram_width = 36;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 11;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 2047;
defparam ram_block1a25.port_a_logical_ram_depth = 2048;
defparam ram_block1a25.port_a_logical_ram_width = 36;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 11;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 2047;
defparam ram_block1a25.port_b_logical_ram_depth = 2048;
defparam ram_block1a25.port_b_logical_ram_width = 36;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 11;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 2047;
defparam ram_block1a30.port_a_logical_ram_depth = 2048;
defparam ram_block1a30.port_a_logical_ram_width = 36;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 11;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 2047;
defparam ram_block1a30.port_b_logical_ram_depth = 2048;
defparam ram_block1a30.port_b_logical_ram_width = 36;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 11;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 2047;
defparam ram_block1a26.port_a_logical_ram_depth = 2048;
defparam ram_block1a26.port_a_logical_ram_width = 36;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 11;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 2047;
defparam ram_block1a26.port_b_logical_ram_depth = 2048;
defparam ram_block1a26.port_b_logical_ram_width = 36;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 11;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 2047;
defparam ram_block1a31.port_a_logical_ram_depth = 2048;
defparam ram_block1a31.port_a_logical_ram_width = 36;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 11;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 2047;
defparam ram_block1a31.port_b_logical_ram_depth = 2048;
defparam ram_block1a31.port_b_logical_ram_width = 36;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 11;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 2047;
defparam ram_block1a27.port_a_logical_ram_depth = 2048;
defparam ram_block1a27.port_a_logical_ram_width = 36;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 11;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 2047;
defparam ram_block1a27.port_b_logical_ram_depth = 2048;
defparam ram_block1a27.port_b_logical_ram_width = 36;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 11;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 2047;
defparam ram_block1a20.port_a_logical_ram_depth = 2048;
defparam ram_block1a20.port_a_logical_ram_width = 36;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 11;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 2047;
defparam ram_block1a20.port_b_logical_ram_depth = 2048;
defparam ram_block1a20.port_b_logical_ram_width = 36;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 11;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 2047;
defparam ram_block1a16.port_a_logical_ram_depth = 2048;
defparam ram_block1a16.port_a_logical_ram_width = 36;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 11;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 2047;
defparam ram_block1a16.port_b_logical_ram_depth = 2048;
defparam ram_block1a16.port_b_logical_ram_width = 36;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 11;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 2047;
defparam ram_block1a21.port_a_logical_ram_depth = 2048;
defparam ram_block1a21.port_a_logical_ram_width = 36;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 11;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 2047;
defparam ram_block1a21.port_b_logical_ram_depth = 2048;
defparam ram_block1a21.port_b_logical_ram_width = 36;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 11;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 2047;
defparam ram_block1a17.port_a_logical_ram_depth = 2048;
defparam ram_block1a17.port_a_logical_ram_width = 36;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 11;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 2047;
defparam ram_block1a17.port_b_logical_ram_depth = 2048;
defparam ram_block1a17.port_b_logical_ram_width = 36;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 11;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 2047;
defparam ram_block1a22.port_a_logical_ram_depth = 2048;
defparam ram_block1a22.port_a_logical_ram_width = 36;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 11;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 2047;
defparam ram_block1a22.port_b_logical_ram_depth = 2048;
defparam ram_block1a22.port_b_logical_ram_width = 36;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 11;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 2047;
defparam ram_block1a18.port_a_logical_ram_depth = 2048;
defparam ram_block1a18.port_a_logical_ram_width = 36;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 11;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 2047;
defparam ram_block1a18.port_b_logical_ram_depth = 2048;
defparam ram_block1a18.port_b_logical_ram_width = 36;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 11;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 2047;
defparam ram_block1a23.port_a_logical_ram_depth = 2048;
defparam ram_block1a23.port_a_logical_ram_width = 36;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 11;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 2047;
defparam ram_block1a23.port_b_logical_ram_depth = 2048;
defparam ram_block1a23.port_b_logical_ram_width = 36;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 11;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 2047;
defparam ram_block1a19.port_a_logical_ram_depth = 2048;
defparam ram_block1a19.port_a_logical_ram_width = 36;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 11;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 2047;
defparam ram_block1a19.port_b_logical_ram_depth = 2048;
defparam ram_block1a19.port_b_logical_ram_width = 36;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 11;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 2047;
defparam ram_block1a12.port_a_logical_ram_depth = 2048;
defparam ram_block1a12.port_a_logical_ram_width = 36;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 11;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 2047;
defparam ram_block1a12.port_b_logical_ram_depth = 2048;
defparam ram_block1a12.port_b_logical_ram_width = 36;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 11;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 2047;
defparam ram_block1a8.port_a_logical_ram_depth = 2048;
defparam ram_block1a8.port_a_logical_ram_width = 36;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 11;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 2047;
defparam ram_block1a8.port_b_logical_ram_depth = 2048;
defparam ram_block1a8.port_b_logical_ram_width = 36;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 11;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 2047;
defparam ram_block1a13.port_a_logical_ram_depth = 2048;
defparam ram_block1a13.port_a_logical_ram_width = 36;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 11;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 2047;
defparam ram_block1a13.port_b_logical_ram_depth = 2048;
defparam ram_block1a13.port_b_logical_ram_width = 36;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 11;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 2047;
defparam ram_block1a9.port_a_logical_ram_depth = 2048;
defparam ram_block1a9.port_a_logical_ram_width = 36;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 11;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 2047;
defparam ram_block1a9.port_b_logical_ram_depth = 2048;
defparam ram_block1a9.port_b_logical_ram_width = 36;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 11;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 2047;
defparam ram_block1a14.port_a_logical_ram_depth = 2048;
defparam ram_block1a14.port_a_logical_ram_width = 36;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 11;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 2047;
defparam ram_block1a14.port_b_logical_ram_depth = 2048;
defparam ram_block1a14.port_b_logical_ram_width = 36;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 11;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 2047;
defparam ram_block1a10.port_a_logical_ram_depth = 2048;
defparam ram_block1a10.port_a_logical_ram_width = 36;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 11;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 2047;
defparam ram_block1a10.port_b_logical_ram_depth = 2048;
defparam ram_block1a10.port_b_logical_ram_width = 36;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 11;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 2047;
defparam ram_block1a15.port_a_logical_ram_depth = 2048;
defparam ram_block1a15.port_a_logical_ram_width = 36;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 11;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 2047;
defparam ram_block1a15.port_b_logical_ram_depth = 2048;
defparam ram_block1a15.port_b_logical_ram_width = 36;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 11;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 2047;
defparam ram_block1a11.port_a_logical_ram_depth = 2048;
defparam ram_block1a11.port_a_logical_ram_width = 36;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 11;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 2047;
defparam ram_block1a11.port_b_logical_ram_depth = 2048;
defparam ram_block1a11.port_b_logical_ram_width = 36;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 11;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 2047;
defparam ram_block1a4.port_a_logical_ram_depth = 2048;
defparam ram_block1a4.port_a_logical_ram_width = 36;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 11;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 2047;
defparam ram_block1a4.port_b_logical_ram_depth = 2048;
defparam ram_block1a4.port_b_logical_ram_width = 36;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 11;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 2047;
defparam ram_block1a0.port_a_logical_ram_depth = 2048;
defparam ram_block1a0.port_a_logical_ram_width = 36;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 11;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 2047;
defparam ram_block1a0.port_b_logical_ram_depth = 2048;
defparam ram_block1a0.port_b_logical_ram_width = 36;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 11;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 2047;
defparam ram_block1a5.port_a_logical_ram_depth = 2048;
defparam ram_block1a5.port_a_logical_ram_width = 36;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 11;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 2047;
defparam ram_block1a5.port_b_logical_ram_depth = 2048;
defparam ram_block1a5.port_b_logical_ram_width = 36;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 11;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 2047;
defparam ram_block1a1.port_a_logical_ram_depth = 2048;
defparam ram_block1a1.port_a_logical_ram_width = 36;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 11;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 2047;
defparam ram_block1a1.port_b_logical_ram_depth = 2048;
defparam ram_block1a1.port_b_logical_ram_width = 36;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 11;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 2047;
defparam ram_block1a6.port_a_logical_ram_depth = 2048;
defparam ram_block1a6.port_a_logical_ram_width = 36;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 11;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 2047;
defparam ram_block1a6.port_b_logical_ram_depth = 2048;
defparam ram_block1a6.port_b_logical_ram_width = 36;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 11;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 2047;
defparam ram_block1a2.port_a_logical_ram_depth = 2048;
defparam ram_block1a2.port_a_logical_ram_width = 36;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 11;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 2047;
defparam ram_block1a2.port_b_logical_ram_depth = 2048;
defparam ram_block1a2.port_b_logical_ram_width = 36;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 11;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 2047;
defparam ram_block1a7.port_a_logical_ram_depth = 2048;
defparam ram_block1a7.port_a_logical_ram_width = 36;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 11;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 2047;
defparam ram_block1a7.port_b_logical_ram_depth = 2048;
defparam ram_block1a7.port_b_logical_ram_width = 36;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(gnd),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_a_fifo_opt_1246:TX_DATA|altera_tse_altsyncram_dpm_fifo:U_RAM|altsyncram:altsyncram_component|altsyncram_3ao1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 11;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 2047;
defparam ram_block1a3.port_a_logical_ram_depth = 2048;
defparam ram_block1a3.port_a_logical_ram_width = 36;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 11;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 2047;
defparam ram_block1a3.port_b_logical_ram_depth = 2048;
defparam ram_block1a3.port_b_logical_ram_width = 36;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_7 (
	reset,
	b_out_10,
	b_out_7,
	b_out_6,
	b_out_3,
	b_out_2,
	b_out_1,
	b_out_0,
	b_out_5,
	b_out_4,
	b_out_9,
	b_out_8,
	always5,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	b_out_10;
output 	b_out_7;
output 	b_out_6;
output 	b_out_3;
output 	b_out_2;
output 	b_out_1;
output 	b_out_0;
output 	b_out_5;
output 	b_out_4;
output 	b_out_9;
output 	b_out_8;
input 	always5;
output 	g_out_10;
output 	g_out_9;
output 	g_out_8;
output 	g_out_7;
output 	g_out_6;
output 	g_out_5;
output 	g_out_4;
output 	g_out_3;
output 	g_out_2;
output 	g_out_1;
output 	g_out_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~25_sumout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \LessThan0~2_combout ;
wire \b_int~0_combout ;
wire \b_int[0]~q ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \b_int[1]~q ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \b_int[2]~q ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \b_int[3]~q ;
wire \Add0~14 ;
wire \Add0~33_sumout ;
wire \b_int[4]~q ;
wire \Add0~34 ;
wire \Add0~29_sumout ;
wire \b_int[5]~q ;
wire \Add0~30 ;
wire \Add0~9_sumout ;
wire \b_int[6]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \b_int[7]~q ;
wire \Add0~6 ;
wire \Add0~41_sumout ;
wire \b_int[8]~q ;
wire \Add0~42 ;
wire \Add0~37_sumout ;
wire \b_int[9]~q ;
wire \Add0~38 ;
wire \Add0~1_sumout ;
wire \b_int[10]~q ;
wire \b_out[0]~0_combout ;
wire \gry_grayval[9]~combout ;
wire \gry_grayval[8]~combout ;
wire \gry_grayval[7]~combout ;
wire \gry_grayval[6]~combout ;
wire \gry_grayval[5]~combout ;
wire \gry_grayval[4]~combout ;
wire \gry_grayval[3]~combout ;
wire \gry_grayval[2]~combout ;
wire \gry_grayval[1]~combout ;
wire \gry_grayval[0]~combout ;


dffeas \b_out[10] (
	.clk(clk),
	.d(\b_int[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_10),
	.prn(vcc));
defparam \b_out[10] .is_wysiwyg = "true";
defparam \b_out[10] .power_up = "low";

dffeas \b_out[7] (
	.clk(clk),
	.d(\b_int[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[6] (
	.clk(clk),
	.d(\b_int[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[3] (
	.clk(clk),
	.d(\b_int[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[2] (
	.clk(clk),
	.d(\b_int[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[1] (
	.clk(clk),
	.d(\b_int[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[0] (
	.clk(clk),
	.d(\b_out[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[5] (
	.clk(clk),
	.d(\b_int[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[4] (
	.clk(clk),
	.d(\b_int[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[9] (
	.clk(clk),
	.d(\b_int[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_9),
	.prn(vcc));
defparam \b_out[9] .is_wysiwyg = "true";
defparam \b_out[9] .power_up = "low";

dffeas \b_out[8] (
	.clk(clk),
	.d(\b_int[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

dffeas \g_out[10] (
	.clk(clk),
	.d(\b_int[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_10),
	.prn(vcc));
defparam \g_out[10] .is_wysiwyg = "true";
defparam \g_out[10] .power_up = "low";

dffeas \g_out[9] (
	.clk(clk),
	.d(\gry_grayval[9]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_9),
	.prn(vcc));
defparam \g_out[9] .is_wysiwyg = "true";
defparam \g_out[9] .power_up = "low";

dffeas \g_out[8] (
	.clk(clk),
	.d(\gry_grayval[8]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_8),
	.prn(vcc));
defparam \g_out[8] .is_wysiwyg = "true";
defparam \g_out[8] .power_up = "low";

dffeas \g_out[7] (
	.clk(clk),
	.d(\gry_grayval[7]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_7),
	.prn(vcc));
defparam \g_out[7] .is_wysiwyg = "true";
defparam \g_out[7] .power_up = "low";

dffeas \g_out[6] (
	.clk(clk),
	.d(\gry_grayval[6]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_6),
	.prn(vcc));
defparam \g_out[6] .is_wysiwyg = "true";
defparam \g_out[6] .power_up = "low";

dffeas \g_out[5] (
	.clk(clk),
	.d(\gry_grayval[5]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_5),
	.prn(vcc));
defparam \g_out[5] .is_wysiwyg = "true";
defparam \g_out[5] .power_up = "low";

dffeas \g_out[4] (
	.clk(clk),
	.d(\gry_grayval[4]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[3] (
	.clk(clk),
	.d(\gry_grayval[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[2] (
	.clk(clk),
	.d(\gry_grayval[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[1] (
	.clk(clk),
	.d(\gry_grayval[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[0] (
	.clk(clk),
	.d(\gry_grayval[0]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\b_int[10]~q ),
	.datab(!\b_int[9]~q ),
	.datac(!\b_int[8]~q ),
	.datad(!\b_int[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\b_int[6]~q ),
	.datab(!\b_int[4]~q ),
	.datac(!\b_int[3]~q ),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~2 (
	.dataa(!\b_int[7]~q ),
	.datab(!\b_int[5]~q ),
	.datac(!\b_int[1]~q ),
	.datad(!\LessThan0~0_combout ),
	.datae(!\LessThan0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~2 .extended_lut = "off";
defparam \LessThan0~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan0~2 .shared_arith = "off";

cyclonev_lcell_comb \b_int~0 (
	.dataa(!\Add0~25_sumout ),
	.datab(!\LessThan0~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_int~0 .extended_lut = "off";
defparam \b_int~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \b_int~0 .shared_arith = "off";

dffeas \b_int[0] (
	.clk(clk),
	.d(\b_int~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[0]~q ),
	.prn(vcc));
defparam \b_int[0] .is_wysiwyg = "true";
defparam \b_int[0] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \b_int[1] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[1]~q ),
	.prn(vcc));
defparam \b_int[1] .is_wysiwyg = "true";
defparam \b_int[1] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \b_int[2] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[2]~q ),
	.prn(vcc));
defparam \b_int[2] .is_wysiwyg = "true";
defparam \b_int[2] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \b_int[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[3]~q ),
	.prn(vcc));
defparam \b_int[3] .is_wysiwyg = "true";
defparam \b_int[3] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \b_int[4] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[4]~q ),
	.prn(vcc));
defparam \b_int[4] .is_wysiwyg = "true";
defparam \b_int[4] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \b_int[5] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[5]~q ),
	.prn(vcc));
defparam \b_int[5] .is_wysiwyg = "true";
defparam \b_int[5] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \b_int[6] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[6]~q ),
	.prn(vcc));
defparam \b_int[6] .is_wysiwyg = "true";
defparam \b_int[6] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \b_int[7] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[7]~q ),
	.prn(vcc));
defparam \b_int[7] .is_wysiwyg = "true";
defparam \b_int[7] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \b_int[8] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[8]~q ),
	.prn(vcc));
defparam \b_int[8] .is_wysiwyg = "true";
defparam \b_int[8] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \b_int[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[9]~q ),
	.prn(vcc));
defparam \b_int[9] .is_wysiwyg = "true";
defparam \b_int[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\b_int[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \b_int[10] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(\LessThan0~2_combout ),
	.sload(gnd),
	.ena(always5),
	.q(\b_int[10]~q ),
	.prn(vcc));
defparam \b_int[10] .is_wysiwyg = "true";
defparam \b_int[10] .power_up = "low";

cyclonev_lcell_comb \b_out[0]~0 (
	.dataa(!\b_int[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[0]~0 .extended_lut = "off";
defparam \b_out[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \b_out[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[9] (
	.dataa(!\b_int[10]~q ),
	.datab(!\b_int[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[9] .extended_lut = "off";
defparam \gry_grayval[9] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[9] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[8] (
	.dataa(!\b_int[9]~q ),
	.datab(!\b_int[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[8] .extended_lut = "off";
defparam \gry_grayval[8] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[8] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[7] (
	.dataa(!\b_int[8]~q ),
	.datab(!\b_int[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[7] .extended_lut = "off";
defparam \gry_grayval[7] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[7] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[6] (
	.dataa(!\b_int[7]~q ),
	.datab(!\b_int[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[6] .extended_lut = "off";
defparam \gry_grayval[6] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[6] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[5] (
	.dataa(!\b_int[6]~q ),
	.datab(!\b_int[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[5] .extended_lut = "off";
defparam \gry_grayval[5] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[5] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[4] (
	.dataa(!\b_int[5]~q ),
	.datab(!\b_int[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[4] .extended_lut = "off";
defparam \gry_grayval[4] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[4] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[3] (
	.dataa(!\b_int[4]~q ),
	.datab(!\b_int[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[3] .extended_lut = "off";
defparam \gry_grayval[3] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[3] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[2] (
	.dataa(!\b_int[3]~q ),
	.datab(!\b_int[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[2] .extended_lut = "off";
defparam \gry_grayval[2] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[2] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[1] (
	.dataa(!\b_int[2]~q ),
	.datab(!\b_int[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[1] .extended_lut = "off";
defparam \gry_grayval[1] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[1] .shared_arith = "off";

cyclonev_lcell_comb \gry_grayval[0] (
	.dataa(!\b_int[1]~q ),
	.datab(!\b_int[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\gry_grayval[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \gry_grayval[0] .extended_lut = "off";
defparam \gry_grayval[0] .lut_mask = 64'h6666666666666666;
defparam \gry_grayval[0] .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_gray_cnt_8 (
	altera_tse_reset_synchronizer_chain_out,
	b_out_10,
	b_out_1,
	b_out_0,
	b_out_3,
	b_out_2,
	b_out_5,
	b_out_4,
	b_out_7,
	b_out_6,
	b_out_9,
	b_out_8,
	g_out_10,
	g_out_9,
	g_out_8,
	g_out_7,
	g_out_6,
	g_out_5,
	g_out_4,
	g_out_3,
	g_out_2,
	g_out_1,
	g_out_0)/* synthesis synthesis_greybox=1 */;
input 	altera_tse_reset_synchronizer_chain_out;
output 	b_out_10;
output 	b_out_1;
output 	b_out_0;
output 	b_out_3;
output 	b_out_2;
output 	b_out_5;
output 	b_out_4;
output 	b_out_7;
output 	b_out_6;
output 	b_out_9;
output 	b_out_8;
output 	g_out_10;
output 	g_out_9;
output 	g_out_8;
output 	g_out_7;
output 	g_out_6;
output 	g_out_5;
output 	g_out_4;
output 	g_out_3;
output 	g_out_2;
output 	g_out_1;
output 	g_out_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \b_out[10]~0_combout ;
wire \b_out[1]~1_combout ;
wire \b_out[3]~2_combout ;
wire \b_out[2]~3_combout ;
wire \b_out[5]~4_combout ;
wire \b_out[4]~5_combout ;
wire \b_out[7]~6_combout ;
wire \b_out[6]~7_combout ;
wire \b_out[9]~8_combout ;
wire \b_out[8]~9_combout ;
wire \g_out[10]~0_combout ;
wire \g_out[9]~1_combout ;
wire \g_out[8]~2_combout ;
wire \g_out[7]~3_combout ;
wire \g_out[6]~4_combout ;
wire \g_out[5]~5_combout ;
wire \g_out[4]~6_combout ;
wire \g_out[3]~7_combout ;
wire \g_out[2]~8_combout ;
wire \g_out[1]~9_combout ;


dffeas \b_out[10] (
	.clk(gnd),
	.d(\b_out[10]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_10),
	.prn(vcc));
defparam \b_out[10] .is_wysiwyg = "true";
defparam \b_out[10] .power_up = "low";

dffeas \b_out[1] (
	.clk(gnd),
	.d(\b_out[1]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_1),
	.prn(vcc));
defparam \b_out[1] .is_wysiwyg = "true";
defparam \b_out[1] .power_up = "low";

dffeas \b_out[0] (
	.clk(gnd),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_0),
	.prn(vcc));
defparam \b_out[0] .is_wysiwyg = "true";
defparam \b_out[0] .power_up = "low";

dffeas \b_out[3] (
	.clk(gnd),
	.d(\b_out[3]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_3),
	.prn(vcc));
defparam \b_out[3] .is_wysiwyg = "true";
defparam \b_out[3] .power_up = "low";

dffeas \b_out[2] (
	.clk(gnd),
	.d(\b_out[2]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_2),
	.prn(vcc));
defparam \b_out[2] .is_wysiwyg = "true";
defparam \b_out[2] .power_up = "low";

dffeas \b_out[5] (
	.clk(gnd),
	.d(\b_out[5]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_5),
	.prn(vcc));
defparam \b_out[5] .is_wysiwyg = "true";
defparam \b_out[5] .power_up = "low";

dffeas \b_out[4] (
	.clk(gnd),
	.d(\b_out[4]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_4),
	.prn(vcc));
defparam \b_out[4] .is_wysiwyg = "true";
defparam \b_out[4] .power_up = "low";

dffeas \b_out[7] (
	.clk(gnd),
	.d(\b_out[7]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_7),
	.prn(vcc));
defparam \b_out[7] .is_wysiwyg = "true";
defparam \b_out[7] .power_up = "low";

dffeas \b_out[6] (
	.clk(gnd),
	.d(\b_out[6]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_6),
	.prn(vcc));
defparam \b_out[6] .is_wysiwyg = "true";
defparam \b_out[6] .power_up = "low";

dffeas \b_out[9] (
	.clk(gnd),
	.d(\b_out[9]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_9),
	.prn(vcc));
defparam \b_out[9] .is_wysiwyg = "true";
defparam \b_out[9] .power_up = "low";

dffeas \b_out[8] (
	.clk(gnd),
	.d(\b_out[8]~9_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_out_8),
	.prn(vcc));
defparam \b_out[8] .is_wysiwyg = "true";
defparam \b_out[8] .power_up = "low";

dffeas \g_out[10] (
	.clk(gnd),
	.d(\g_out[10]~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_10),
	.prn(vcc));
defparam \g_out[10] .is_wysiwyg = "true";
defparam \g_out[10] .power_up = "low";

dffeas \g_out[9] (
	.clk(gnd),
	.d(\g_out[9]~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_9),
	.prn(vcc));
defparam \g_out[9] .is_wysiwyg = "true";
defparam \g_out[9] .power_up = "low";

dffeas \g_out[8] (
	.clk(gnd),
	.d(\g_out[8]~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_8),
	.prn(vcc));
defparam \g_out[8] .is_wysiwyg = "true";
defparam \g_out[8] .power_up = "low";

dffeas \g_out[7] (
	.clk(gnd),
	.d(\g_out[7]~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_7),
	.prn(vcc));
defparam \g_out[7] .is_wysiwyg = "true";
defparam \g_out[7] .power_up = "low";

dffeas \g_out[6] (
	.clk(gnd),
	.d(\g_out[6]~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_6),
	.prn(vcc));
defparam \g_out[6] .is_wysiwyg = "true";
defparam \g_out[6] .power_up = "low";

dffeas \g_out[5] (
	.clk(gnd),
	.d(\g_out[5]~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_5),
	.prn(vcc));
defparam \g_out[5] .is_wysiwyg = "true";
defparam \g_out[5] .power_up = "low";

dffeas \g_out[4] (
	.clk(gnd),
	.d(\g_out[4]~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_4),
	.prn(vcc));
defparam \g_out[4] .is_wysiwyg = "true";
defparam \g_out[4] .power_up = "low";

dffeas \g_out[3] (
	.clk(gnd),
	.d(\g_out[3]~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_3),
	.prn(vcc));
defparam \g_out[3] .is_wysiwyg = "true";
defparam \g_out[3] .power_up = "low";

dffeas \g_out[2] (
	.clk(gnd),
	.d(\g_out[2]~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_2),
	.prn(vcc));
defparam \g_out[2] .is_wysiwyg = "true";
defparam \g_out[2] .power_up = "low";

dffeas \g_out[1] (
	.clk(gnd),
	.d(\g_out[1]~9_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_1),
	.prn(vcc));
defparam \g_out[1] .is_wysiwyg = "true";
defparam \g_out[1] .power_up = "low";

dffeas \g_out[0] (
	.clk(gnd),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(g_out_0),
	.prn(vcc));
defparam \g_out[0] .is_wysiwyg = "true";
defparam \g_out[0] .power_up = "low";

cyclonev_lcell_comb \b_out[10]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[10]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[10]~0 .extended_lut = "off";
defparam \b_out[10]~0 .lut_mask = 64'h0000000000000000;
defparam \b_out[10]~0 .shared_arith = "off";

cyclonev_lcell_comb \b_out[1]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[1]~1 .extended_lut = "off";
defparam \b_out[1]~1 .lut_mask = 64'h0000000000000000;
defparam \b_out[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \b_out[3]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[3]~2 .extended_lut = "off";
defparam \b_out[3]~2 .lut_mask = 64'h0000000000000000;
defparam \b_out[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \b_out[2]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[2]~3 .extended_lut = "off";
defparam \b_out[2]~3 .lut_mask = 64'h0000000000000000;
defparam \b_out[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \b_out[5]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[5]~4 .extended_lut = "off";
defparam \b_out[5]~4 .lut_mask = 64'h0000000000000000;
defparam \b_out[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \b_out[4]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[4]~5 .extended_lut = "off";
defparam \b_out[4]~5 .lut_mask = 64'h0000000000000000;
defparam \b_out[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \b_out[7]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[7]~6 .extended_lut = "off";
defparam \b_out[7]~6 .lut_mask = 64'h0000000000000000;
defparam \b_out[7]~6 .shared_arith = "off";

cyclonev_lcell_comb \b_out[6]~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[6]~7 .extended_lut = "off";
defparam \b_out[6]~7 .lut_mask = 64'h0000000000000000;
defparam \b_out[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \b_out[9]~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[9]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[9]~8 .extended_lut = "off";
defparam \b_out[9]~8 .lut_mask = 64'h0000000000000000;
defparam \b_out[9]~8 .shared_arith = "off";

cyclonev_lcell_comb \b_out[8]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_out[8]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_out[8]~9 .extended_lut = "off";
defparam \b_out[8]~9 .lut_mask = 64'h0000000000000000;
defparam \b_out[8]~9 .shared_arith = "off";

cyclonev_lcell_comb \g_out[10]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[10]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[10]~0 .extended_lut = "off";
defparam \g_out[10]~0 .lut_mask = 64'h0000000000000000;
defparam \g_out[10]~0 .shared_arith = "off";

cyclonev_lcell_comb \g_out[9]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[9]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[9]~1 .extended_lut = "off";
defparam \g_out[9]~1 .lut_mask = 64'h0000000000000000;
defparam \g_out[9]~1 .shared_arith = "off";

cyclonev_lcell_comb \g_out[8]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[8]~2 .extended_lut = "off";
defparam \g_out[8]~2 .lut_mask = 64'h0000000000000000;
defparam \g_out[8]~2 .shared_arith = "off";

cyclonev_lcell_comb \g_out[7]~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[7]~3 .extended_lut = "off";
defparam \g_out[7]~3 .lut_mask = 64'h0000000000000000;
defparam \g_out[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \g_out[6]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[6]~4 .extended_lut = "off";
defparam \g_out[6]~4 .lut_mask = 64'h0000000000000000;
defparam \g_out[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \g_out[5]~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[5]~5 .extended_lut = "off";
defparam \g_out[5]~5 .lut_mask = 64'h0000000000000000;
defparam \g_out[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \g_out[4]~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[4]~6 .extended_lut = "off";
defparam \g_out[4]~6 .lut_mask = 64'h0000000000000000;
defparam \g_out[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \g_out[3]~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[3]~7 .extended_lut = "off";
defparam \g_out[3]~7 .lut_mask = 64'h0000000000000000;
defparam \g_out[3]~7 .shared_arith = "off";

cyclonev_lcell_comb \g_out[2]~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[2]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[2]~8 .extended_lut = "off";
defparam \g_out[2]~8 .lut_mask = 64'h0000000000000000;
defparam \g_out[2]~8 .shared_arith = "off";

cyclonev_lcell_comb \g_out[1]~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\g_out[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \g_out[1]~9 .extended_lut = "off";
defparam \g_out[1]~9 .lut_mask = 64'h0000000000000000;
defparam \g_out[1]~9 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_altsyncram_dpm_fifo_4 (
	q_b_9,
	eop_sft_0,
	transmit_cnt_0,
	transmit_cnt_1,
	transmit_cnt_2,
	transmit_cnt_3,
	transmit_cnt_4,
	transmit_cnt_5,
	transmit_cnt_6,
	q_b_8,
	q_b_4,
	dout_reg_sft_28,
	q_b_0,
	dout_reg_sft_24,
	q_b_5,
	dout_reg_sft_29,
	q_b_1,
	dout_reg_sft_25,
	q_b_6,
	dout_reg_sft_30,
	q_b_2,
	dout_reg_sft_26,
	q_b_7,
	dout_reg_sft_31,
	q_b_3,
	dout_reg_sft_27,
	buf_wren,
	buf_wraddr_0,
	buf_wraddr_1,
	buf_wraddr_2,
	buf_wraddr_3,
	buf_wraddr_4,
	buf_wraddr_5,
	buf_wraddr_6,
	sop_reg,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_9;
input 	eop_sft_0;
input 	transmit_cnt_0;
input 	transmit_cnt_1;
input 	transmit_cnt_2;
input 	transmit_cnt_3;
input 	transmit_cnt_4;
input 	transmit_cnt_5;
input 	transmit_cnt_6;
output 	q_b_8;
output 	q_b_4;
input 	dout_reg_sft_28;
output 	q_b_0;
input 	dout_reg_sft_24;
output 	q_b_5;
input 	dout_reg_sft_29;
output 	q_b_1;
input 	dout_reg_sft_25;
output 	q_b_6;
input 	dout_reg_sft_30;
output 	q_b_2;
input 	dout_reg_sft_26;
output 	q_b_7;
input 	dout_reg_sft_31;
output 	q_b_3;
input 	dout_reg_sft_27;
input 	buf_wren;
input 	buf_wraddr_0;
input 	buf_wraddr_1;
input 	buf_wraddr_2;
input 	buf_wraddr_3;
input 	buf_wraddr_4;
input 	buf_wraddr_5;
input 	buf_wraddr_6;
input 	sop_reg;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_6 altsyncram_component(
	.q_b({q_b_unconnected_wire_39,q_b_unconnected_wire_38,q_b_unconnected_wire_37,q_b_unconnected_wire_36,q_b_unconnected_wire_35,q_b_unconnected_wire_34,q_b_unconnected_wire_33,q_b_unconnected_wire_32,q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,
q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,
q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,eop_sft_0,sop_reg,dout_reg_sft_31,dout_reg_sft_30,dout_reg_sft_29,dout_reg_sft_28,dout_reg_sft_27,dout_reg_sft_26,dout_reg_sft_25,dout_reg_sft_24}),
	.address_b({gnd,gnd,gnd,gnd,transmit_cnt_6,transmit_cnt_5,transmit_cnt_4,transmit_cnt_3,transmit_cnt_2,transmit_cnt_1,transmit_cnt_0}),
	.wren_a(buf_wren),
	.address_a({gnd,gnd,gnd,gnd,buf_wraddr_6,buf_wraddr_5,buf_wraddr_4,buf_wraddr_3,buf_wraddr_2,buf_wraddr_1,buf_wraddr_0}),
	.clock0(mac_tx_clock_connection_clk));

endmodule

module IoTOctopus_QSYS_altsyncram_6 (
	q_b,
	data_a,
	address_b,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[39:0] q_b;
input 	[39:0] data_a;
input 	[10:0] address_b;
input 	wren_a;
input 	[10:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



IoTOctopus_QSYS_altsyncram_n3o1 auto_generated(
	.q_b({q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0),
	.clock1(clock0));

endmodule

module IoTOctopus_QSYS_altsyncram_n3o1 (
	q_b,
	data_a,
	address_b,
	wren_a,
	address_a,
	clock0,
	clock1)/* synthesis synthesis_greybox=1 */;
output 	[9:0] q_b;
input 	[9:0] data_a;
input 	[6:0] address_b;
input 	wren_a;
input 	[6:0] address_a;
input 	clock0;
input 	clock1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 10;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 10;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 10;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 10;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 10;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 10;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 10;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 10;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 10;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "IoTOctopus_QSYS_eth_tse_0:eth_tse_0|altera_eth_tse_mac:i_tse_mac|altera_tse_top_w_fifo_10_100_1000:U_MAC_TOP|altera_tse_top_w_fifo:U_MAC|altera_tse_tx_min_ff:U_TXFF|altera_tse_altsyncram_dpm_fifo:U_RTSM|altsyncram:altsyncram_component|altsyncram_n3o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 10;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

endmodule

module IoTOctopus_QSYS_altera_tse_retransmit_cntl (
	q_b_9,
	eop_sft_0,
	transmit_cnt_0,
	transmit_cnt_1,
	transmit_cnt_2,
	transmit_cnt_3,
	transmit_cnt_4,
	transmit_cnt_5,
	transmit_cnt_6,
	clk_ena,
	altera_tse_reset_synchronizer_chain_out,
	dreg_1,
	retrans_ena1,
	dreg_11,
	always9,
	buf_wren1,
	buf_wraddr_0,
	buf_wraddr_1,
	buf_wraddr_2,
	buf_wraddr_3,
	buf_wraddr_4,
	buf_wraddr_5,
	buf_wraddr_6,
	stateSTM_TYP_WAIT_COL_1,
	stateSTM_TYP_RETRANSMIT_SHORT,
	col_int,
	Selector4,
	short_frm1,
	always91,
	tx_rden_mii,
	Selector1,
	Selector5,
	always10,
	tx_rden_int,
	Selector3,
	Selector31,
	always92,
	Selector32,
	mac_ena1,
	crs,
	stat_rden1,
	tx_stat_rden,
	GND_port,
	mac_tx_clock_connection_clk)/* synthesis synthesis_greybox=1 */;
input 	q_b_9;
input 	eop_sft_0;
output 	transmit_cnt_0;
output 	transmit_cnt_1;
output 	transmit_cnt_2;
output 	transmit_cnt_3;
output 	transmit_cnt_4;
output 	transmit_cnt_5;
output 	transmit_cnt_6;
input 	clk_ena;
input 	altera_tse_reset_synchronizer_chain_out;
input 	dreg_1;
output 	retrans_ena1;
input 	dreg_11;
input 	always9;
output 	buf_wren1;
output 	buf_wraddr_0;
output 	buf_wraddr_1;
output 	buf_wraddr_2;
output 	buf_wraddr_3;
output 	buf_wraddr_4;
output 	buf_wraddr_5;
output 	buf_wraddr_6;
output 	stateSTM_TYP_WAIT_COL_1;
output 	stateSTM_TYP_RETRANSMIT_SHORT;
input 	col_int;
output 	Selector4;
output 	short_frm1;
input 	always91;
input 	tx_rden_mii;
output 	Selector1;
output 	Selector5;
output 	always10;
input 	tx_rden_int;
output 	Selector3;
output 	Selector31;
input 	always92;
output 	Selector32;
output 	mac_ena1;
input 	crs;
output 	stat_rden1;
input 	tx_stat_rden;
input 	GND_port;
input 	mac_tx_clock_connection_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \U_LFSR|z_reg[9]~q ;
wire \U_LFSR|z_reg[8]~q ;
wire \U_LFSR|z_reg[7]~q ;
wire \U_LFSR|z_reg[6]~q ;
wire \U_LFSR|z_reg[5]~q ;
wire \U_LFSR|z_reg[4]~q ;
wire \U_LFSR|z_reg[3]~q ;
wire \U_LFSR|z_reg[2]~q ;
wire \U_LFSR|z_reg[1]~q ;
wire \U_LFSR|z_reg[0]~q ;
wire \lfsr_ena~combout ;
wire \Add4~1_sumout ;
wire \state.STM_TYP_IDLE~0_combout ;
wire \state.STM_TYP_IDLE~q ;
wire \Selector1~0_combout ;
wire \Selector4~4_combout ;
wire \Selector4~1_combout ;
wire \state.STM_TYP_RETRANSMIT~q ;
wire \state.STM_TYP_FLUSH~q ;
wire \load_cnt_reg[3]~q ;
wire \load_cnt_reg[2]~q ;
wire \load_cnt_reg[1]~q ;
wire \load_cnt_reg[0]~q ;
wire \Add3~25_sumout ;
wire \load_cnt~8_combout ;
wire \Selector4~3_combout ;
wire \Selector0~7_combout ;
wire \load_cnt_reg[4]~q ;
wire \Add3~14 ;
wire \Add3~9_sumout ;
wire \load_cnt~4_combout ;
wire \load_cnt[4]~q ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \load_cnt[6]~1_combout ;
wire \load_cnt[6]~2_combout ;
wire \load_cnt[0]~q ;
wire \Add3~26 ;
wire \Add3~21_sumout ;
wire \load_cnt~7_combout ;
wire \load_cnt[1]~q ;
wire \Add3~22 ;
wire \Add3~17_sumout ;
wire \load_cnt~6_combout ;
wire \load_cnt[2]~q ;
wire \Add3~18 ;
wire \Add3~13_sumout ;
wire \load_cnt~5_combout ;
wire \load_cnt[3]~q ;
wire \LessThan0~0_combout ;
wire \Selector2~0_combout ;
wire \state.STM_TYP_WAIT_END~q ;
wire \Selector7~5_combout ;
wire \Add1~1_sumout ;
wire \Add2~1_sumout ;
wire \Add0~1_sumout ;
wire \wait_col_cnt~0_combout ;
wire \Equal1~1_combout ;
wire \Equal1~2_combout ;
wire \Selector1~2_combout ;
wire \Selector1~3_combout ;
wire \Add1~2 ;
wire \Add1~26 ;
wire \Add1~22 ;
wire \Add1~18 ;
wire \Add1~14 ;
wire \Add1~10 ;
wire \Add1~5_sumout ;
wire \Add1~9_sumout ;
wire \Add1~13_sumout ;
wire \Add1~17_sumout ;
wire \Add1~21_sumout ;
wire \Add1~25_sumout ;
wire \Add2~2 ;
wire \Add2~25_sumout ;
wire \Add0~2 ;
wire \Add0~25_sumout ;
wire \wait_col_cnt~8_combout ;
wire \wait_col_cnt[1]~q ;
wire \Add2~26 ;
wire \Add2~21_sumout ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \wait_col_cnt~7_combout ;
wire \wait_col_cnt[2]~q ;
wire \Add2~22 ;
wire \Add2~17_sumout ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \wait_col_cnt~6_combout ;
wire \wait_col_cnt[3]~q ;
wire \Add2~18 ;
wire \Add2~13_sumout ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \wait_col_cnt~5_combout ;
wire \wait_col_cnt[4]~q ;
wire \Add2~14 ;
wire \Add2~9_sumout ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \wait_col_cnt~4_combout ;
wire \wait_col_cnt[5]~q ;
wire \Add2~10 ;
wire \Add2~5_sumout ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \wait_col_cnt~3_combout ;
wire \wait_col_cnt[6]~q ;
wire \Equal0~0_combout ;
wire \Selector7~6_combout ;
wire \wait_col_cnt[6]~1_combout ;
wire \wait_col_cnt[6]~2_combout ;
wire \wait_col_cnt[0]~q ;
wire \always0~4_combout ;
wire \Selector7~3_combout ;
wire \Selector7~4_combout ;
wire \state.STM_TYP_WAIT_COL~q ;
wire \Add6~13_sumout ;
wire \always14~0_combout ;
wire \Add6~2 ;
wire \Add6~61_sumout ;
wire \back_cnt[4]~q ;
wire \Add6~62 ;
wire \Add6~57_sumout ;
wire \back_cnt[5]~q ;
wire \Add6~58 ;
wire \Add6~53_sumout ;
wire \back_cnt[6]~q ;
wire \Add6~54 ;
wire \Add6~49_sumout ;
wire \wait_late~0_combout ;
wire \wait_late~1_combout ;
wire \wait_late~2_combout ;
wire \wait_late~3_combout ;
wire \wait_late~q ;
wire \Selector6~2_combout ;
wire \Selector6~8_combout ;
wire \Selector6~6_combout ;
wire \retrans_cnt~0_combout ;
wire \retrans_cnt~7_combout ;
wire \retrans_cnt[3]~2_combout ;
wire \retrans_cnt[3]~3_combout ;
wire \retrans_cnt[0]~q ;
wire \Add5~3_combout ;
wire \retrans_cnt~6_combout ;
wire \retrans_cnt[1]~q ;
wire \Add5~2_combout ;
wire \retrans_cnt~5_combout ;
wire \retrans_cnt[2]~q ;
wire \Add5~1_combout ;
wire \retrans_cnt~4_combout ;
wire \retrans_cnt[3]~q ;
wire \Equal3~0_combout ;
wire \back_cnt~9_combout ;
wire \back_cnt[7]~q ;
wire \Add6~50 ;
wire \Add6~45_sumout ;
wire \back_cnt~8_combout ;
wire \back_cnt[8]~q ;
wire \Add6~46 ;
wire \Add6~41_sumout ;
wire \back_cnt~7_combout ;
wire \back_cnt[9]~q ;
wire \Add6~42 ;
wire \Add6~37_sumout ;
wire \back_cnt~6_combout ;
wire \back_cnt[10]~q ;
wire \Add6~38 ;
wire \Add6~33_sumout ;
wire \back_cnt~5_combout ;
wire \back_cnt[11]~q ;
wire \Add6~34 ;
wire \Add6~29_sumout ;
wire \back_cnt~4_combout ;
wire \back_cnt[12]~q ;
wire \Add6~30 ;
wire \Add6~25_sumout ;
wire \back_cnt~3_combout ;
wire \back_cnt[13]~q ;
wire \Add6~26 ;
wire \Add6~21_sumout ;
wire \back_cnt~2_combout ;
wire \back_cnt[14]~q ;
wire \Add6~22 ;
wire \Add6~17_sumout ;
wire \back_cnt~1_combout ;
wire \back_cnt[15]~q ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \Equal2~3_combout ;
wire \Selector6~7_combout ;
wire \Selector6~5_combout ;
wire \back_cnt~0_combout ;
wire \back_cnt[0]~q ;
wire \Add6~14 ;
wire \Add6~9_sumout ;
wire \back_cnt[1]~q ;
wire \Add6~10 ;
wire \Add6~5_sumout ;
wire \back_cnt[2]~q ;
wire \Add6~6 ;
wire \Add6~1_sumout ;
wire \back_cnt[3]~q ;
wire \Equal2~0_combout ;
wire \Selector6~1_combout ;
wire \Add5~0_combout ;
wire \retrans_cnt~1_combout ;
wire \retrans_cnt[4]~q ;
wire \always16~0_combout ;
wire \excess_col_int~q ;
wire \Selector0~2_combout ;
wire \col_reg~0_combout ;
wire \col_reg~q ;
wire \Selector1~4_combout ;
wire \state.STM_TYP_COPY~q ;
wire \load_cnt_reg~0_combout ;
wire \load_cnt_reg[5]~q ;
wire \Add3~10 ;
wire \Add3~5_sumout ;
wire \load_cnt~3_combout ;
wire \load_cnt[5]~q ;
wire \Add3~6 ;
wire \Add3~1_sumout ;
wire \load_cnt~0_combout ;
wire \load_cnt[6]~q ;
wire \load_cnt_reg[6]~q ;
wire \Equal1~0_combout ;
wire \Selector4~2_combout ;
wire \Selector6~3_combout ;
wire \Selector6~4_combout ;
wire \state.STM_TYP_BACK_OFF~q ;
wire \Selector0~3_combout ;
wire \Selector0~4_combout ;
wire \Selector0~5_combout ;
wire \Selector0~8_combout ;
wire \Selector0~6_combout ;
wire \Selector5~1_combout ;
wire \Selector5~3_combout ;
wire \Selector5~2_combout ;
wire \clk_ena_reg~q ;
wire \mac_ff_rden_reg~0_combout ;
wire \mac_ff_rden_reg~q ;
wire \transmit_cnt[6]~0_combout ;
wire \Add4~2 ;
wire \Add4~5_sumout ;
wire \Add4~6 ;
wire \Add4~9_sumout ;
wire \Add4~10 ;
wire \Add4~13_sumout ;
wire \Add4~14 ;
wire \Add4~17_sumout ;
wire \Add4~18 ;
wire \Add4~21_sumout ;
wire \Add4~22 ;
wire \Add4~25_sumout ;
wire \always9~0_combout ;
wire \Selector8~0_combout ;
wire \always0~3_combout ;
wire \always0~5_combout ;
wire \short_frm~0_combout ;
wire \always10~1_combout ;
wire \always10~2_combout ;
wire \Selector3~1_combout ;
wire \crs_d~q ;
wire \mac_ena~0_combout ;
wire \mac_ena~1_combout ;
wire \mac_ena~2_combout ;
wire \mac_ena~3_combout ;
wire \stat_rden~0_combout ;


IoTOctopus_QSYS_altera_tse_lfsr_10 U_LFSR(
	.reset(altera_tse_reset_synchronizer_chain_out),
	.z_reg_9(\U_LFSR|z_reg[9]~q ),
	.z_reg_8(\U_LFSR|z_reg[8]~q ),
	.z_reg_7(\U_LFSR|z_reg[7]~q ),
	.z_reg_6(\U_LFSR|z_reg[6]~q ),
	.z_reg_5(\U_LFSR|z_reg[5]~q ),
	.z_reg_4(\U_LFSR|z_reg[4]~q ),
	.z_reg_3(\U_LFSR|z_reg[3]~q ),
	.z_reg_2(\U_LFSR|z_reg[2]~q ),
	.z_reg_1(\U_LFSR|z_reg[1]~q ),
	.z_reg_0(\U_LFSR|z_reg[0]~q ),
	.enable(\lfsr_ena~combout ),
	.tx_clk(mac_tx_clock_connection_clk));

cyclonev_lcell_comb lfsr_ena(
	.dataa(!clk_ena),
	.datab(!dreg_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_ena~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam lfsr_ena.extended_lut = "off";
defparam lfsr_ena.lut_mask = 64'h7777777777777777;
defparam lfsr_ena.shared_arith = "off";

dffeas \transmit_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~1_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_0),
	.prn(vcc));
defparam \transmit_cnt[0] .is_wysiwyg = "true";
defparam \transmit_cnt[0] .power_up = "low";

dffeas \transmit_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~5_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_1),
	.prn(vcc));
defparam \transmit_cnt[1] .is_wysiwyg = "true";
defparam \transmit_cnt[1] .power_up = "low";

dffeas \transmit_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~9_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_2),
	.prn(vcc));
defparam \transmit_cnt[2] .is_wysiwyg = "true";
defparam \transmit_cnt[2] .power_up = "low";

dffeas \transmit_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~13_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_3),
	.prn(vcc));
defparam \transmit_cnt[3] .is_wysiwyg = "true";
defparam \transmit_cnt[3] .power_up = "low";

dffeas \transmit_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~17_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_4),
	.prn(vcc));
defparam \transmit_cnt[4] .is_wysiwyg = "true";
defparam \transmit_cnt[4] .power_up = "low";

dffeas \transmit_cnt[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~21_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_5),
	.prn(vcc));
defparam \transmit_cnt[5] .is_wysiwyg = "true";
defparam \transmit_cnt[5] .power_up = "low";

dffeas \transmit_cnt[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add4~25_sumout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\transmit_cnt[6]~0_combout ),
	.q(transmit_cnt_6),
	.prn(vcc));
defparam \transmit_cnt[6] .is_wysiwyg = "true";
defparam \transmit_cnt[6] .power_up = "low";

dffeas retrans_ena(
	.clk(mac_tx_clock_connection_clk),
	.d(always10),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(retrans_ena1),
	.prn(vcc));
defparam retrans_ena.is_wysiwyg = "true";
defparam retrans_ena.power_up = "low";

dffeas buf_wren(
	.clk(mac_tx_clock_connection_clk),
	.d(\always9~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wren1),
	.prn(vcc));
defparam buf_wren.is_wysiwyg = "true";
defparam buf_wren.power_up = "low";

dffeas \buf_wraddr[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_0),
	.prn(vcc));
defparam \buf_wraddr[0] .is_wysiwyg = "true";
defparam \buf_wraddr[0] .power_up = "low";

dffeas \buf_wraddr[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_1),
	.prn(vcc));
defparam \buf_wraddr[1] .is_wysiwyg = "true";
defparam \buf_wraddr[1] .power_up = "low";

dffeas \buf_wraddr[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_2),
	.prn(vcc));
defparam \buf_wraddr[2] .is_wysiwyg = "true";
defparam \buf_wraddr[2] .power_up = "low";

dffeas \buf_wraddr[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_3),
	.prn(vcc));
defparam \buf_wraddr[3] .is_wysiwyg = "true";
defparam \buf_wraddr[3] .power_up = "low";

dffeas \buf_wraddr[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_4),
	.prn(vcc));
defparam \buf_wraddr[4] .is_wysiwyg = "true";
defparam \buf_wraddr[4] .power_up = "low";

dffeas \buf_wraddr[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_5),
	.prn(vcc));
defparam \buf_wraddr[5] .is_wysiwyg = "true";
defparam \buf_wraddr[5] .power_up = "low";

dffeas \buf_wraddr[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(buf_wraddr_6),
	.prn(vcc));
defparam \buf_wraddr[6] .is_wysiwyg = "true";
defparam \buf_wraddr[6] .power_up = "low";

dffeas \state.STM_TYP_WAIT_COL_1 (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateSTM_TYP_WAIT_COL_1),
	.prn(vcc));
defparam \state.STM_TYP_WAIT_COL_1 .is_wysiwyg = "true";
defparam \state.STM_TYP_WAIT_COL_1 .power_up = "low";

dffeas \state.STM_TYP_RETRANSMIT_SHORT (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector5~2_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateSTM_TYP_RETRANSMIT_SHORT),
	.prn(vcc));
defparam \state.STM_TYP_RETRANSMIT_SHORT .is_wysiwyg = "true";
defparam \state.STM_TYP_RETRANSMIT_SHORT .power_up = "low";

cyclonev_lcell_comb \Selector4~0 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_RETRANSMIT~q ),
	.datac(!\Equal1~0_combout ),
	.datad(!\Equal1~1_combout ),
	.datae(!\Equal1~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~0 .extended_lut = "off";
defparam \Selector4~0 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \Selector4~0 .shared_arith = "off";

dffeas short_frm(
	.clk(mac_tx_clock_connection_clk),
	.d(\short_frm~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(short_frm1),
	.prn(vcc));
defparam short_frm.is_wysiwyg = "true";
defparam short_frm.power_up = "low";

cyclonev_lcell_comb \Selector1~1 (
	.dataa(!clk_ena),
	.datab(!dreg_11),
	.datac(!always91),
	.datad(!always9),
	.datae(!tx_rden_mii),
	.dataf(!\Selector1~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~1 .extended_lut = "off";
defparam \Selector1~1 .lut_mask = 64'h47FFFFFFFFFFFFFF;
defparam \Selector1~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~0 (
	.dataa(!dreg_1),
	.datab(!\col_reg~q ),
	.datac(!\excess_col_int~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector5),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~0 .extended_lut = "off";
defparam \Selector5~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Selector5~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~0 (
	.dataa(!\Selector8~0_combout ),
	.datab(!Selector4),
	.datac(!\Selector5~1_combout ),
	.datad(!always91),
	.datae(!\always10~1_combout ),
	.dataf(!\always10~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always10),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~0 .extended_lut = "off";
defparam \always10~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \always10~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~0 (
	.dataa(!dreg_1),
	.datab(!\excess_col_int~q ),
	.datac(!\state.STM_TYP_IDLE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector3),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~0 .extended_lut = "off";
defparam \Selector3~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Selector3~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~2 (
	.dataa(!eop_sft_0),
	.datab(!short_frm1),
	.datac(!\col_reg~q ),
	.datad(!\Selector3~1_combout ),
	.datae(!\state.STM_TYP_FLUSH~q ),
	.dataf(!Selector3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector31),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~2 .extended_lut = "off";
defparam \Selector3~2 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \Selector3~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~3 (
	.dataa(!dreg_11),
	.datab(!always92),
	.datac(!tx_rden_mii),
	.datad(!Selector3),
	.datae(!Selector31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Selector32),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~3 .extended_lut = "off";
defparam \Selector3~3 .lut_mask = 64'hFFFFD8FFFFFFD8FF;
defparam \Selector3~3 .shared_arith = "off";

dffeas mac_ena(
	.clk(mac_tx_clock_connection_clk),
	.d(\mac_ena~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mac_ena1),
	.prn(vcc));
defparam mac_ena.is_wysiwyg = "true";
defparam mac_ena.power_up = "low";

dffeas stat_rden(
	.clk(mac_tx_clock_connection_clk),
	.d(\stat_rden~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stat_rden1),
	.prn(vcc));
defparam stat_rden.is_wysiwyg = "true";
defparam stat_rden.power_up = "low";

cyclonev_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~1_sumout ),
	.cout(\Add4~2 ),
	.shareout());
defparam \Add4~1 .extended_lut = "off";
defparam \Add4~1 .lut_mask = 64'h00000000000000FF;
defparam \Add4~1 .shared_arith = "off";

cyclonev_lcell_comb \state.STM_TYP_IDLE~0 (
	.dataa(!\Selector0~6_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state.STM_TYP_IDLE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state.STM_TYP_IDLE~0 .extended_lut = "off";
defparam \state.STM_TYP_IDLE~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \state.STM_TYP_IDLE~0 .shared_arith = "off";

dffeas \state.STM_TYP_IDLE (
	.clk(mac_tx_clock_connection_clk),
	.d(\state.STM_TYP_IDLE~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_IDLE~q ),
	.prn(vcc));
defparam \state.STM_TYP_IDLE .is_wysiwyg = "true";
defparam \state.STM_TYP_IDLE .power_up = "low";

cyclonev_lcell_comb \Selector1~0 (
	.dataa(!dreg_1),
	.datab(!\state.STM_TYP_IDLE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~0 .extended_lut = "off";
defparam \Selector1~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~4 (
	.dataa(!short_frm1),
	.datab(!clk_ena),
	.datac(!dreg_11),
	.datad(!tx_rden_mii),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~4 .extended_lut = "off";
defparam \Selector4~4 .lut_mask = 64'hA3FFFFFFA3FFFFFF;
defparam \Selector4~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~1 (
	.dataa(!Selector4),
	.datab(!Selector5),
	.datac(!dreg_11),
	.datad(!always91),
	.datae(!always9),
	.dataf(!\Selector4~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~1 .extended_lut = "off";
defparam \Selector4~1 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \Selector4~1 .shared_arith = "off";

dffeas \state.STM_TYP_RETRANSMIT (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector4~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_RETRANSMIT~q ),
	.prn(vcc));
defparam \state.STM_TYP_RETRANSMIT .is_wysiwyg = "true";
defparam \state.STM_TYP_RETRANSMIT .power_up = "low";

dffeas \state.STM_TYP_FLUSH (
	.clk(mac_tx_clock_connection_clk),
	.d(Selector32),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_FLUSH~q ),
	.prn(vcc));
defparam \state.STM_TYP_FLUSH .is_wysiwyg = "true";
defparam \state.STM_TYP_FLUSH .power_up = "low";

dffeas \load_cnt_reg[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[3]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[3]~q ),
	.prn(vcc));
defparam \load_cnt_reg[3] .is_wysiwyg = "true";
defparam \load_cnt_reg[3] .power_up = "low";

dffeas \load_cnt_reg[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[2]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[2]~q ),
	.prn(vcc));
defparam \load_cnt_reg[2] .is_wysiwyg = "true";
defparam \load_cnt_reg[2] .power_up = "low";

dffeas \load_cnt_reg[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[1]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[1]~q ),
	.prn(vcc));
defparam \load_cnt_reg[1] .is_wysiwyg = "true";
defparam \load_cnt_reg[1] .power_up = "low";

dffeas \load_cnt_reg[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[0]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[0]~q ),
	.prn(vcc));
defparam \load_cnt_reg[0] .is_wysiwyg = "true";
defparam \load_cnt_reg[0] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h00000000000000FF;
defparam \Add3~25 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt~8 (
	.dataa(!\load_cnt_reg[0]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~25_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~8 .extended_lut = "off";
defparam \load_cnt~8 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~3 (
	.dataa(!dreg_11),
	.datab(!short_frm1),
	.datac(!always92),
	.datad(!tx_rden_mii),
	.datae(!\Selector1~0_combout ),
	.dataf(!Selector5),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~3 .extended_lut = "off";
defparam \Selector4~3 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \Selector4~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~7 (
	.dataa(!dreg_11),
	.datab(!\excess_col_int~q ),
	.datac(!\state.STM_TYP_IDLE~q ),
	.datad(!always92),
	.datae(!tx_rden_mii),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~7 .extended_lut = "off";
defparam \Selector0~7 .lut_mask = 64'hFFFFFFD8FFFFFFD8;
defparam \Selector0~7 .shared_arith = "off";

dffeas \load_cnt_reg[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[4]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[4]~q ),
	.prn(vcc));
defparam \load_cnt_reg[4] .is_wysiwyg = "true";
defparam \load_cnt_reg[4] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h00000000000000FF;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h00000000000000FF;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt~4 (
	.dataa(!\load_cnt_reg[4]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~4 .extended_lut = "off";
defparam \load_cnt~4 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~4 .shared_arith = "off";

dffeas \load_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[4]~q ),
	.prn(vcc));
defparam \load_cnt[4] .is_wysiwyg = "true";
defparam \load_cnt[4] .power_up = "low";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!\load_cnt[3]~q ),
	.datab(!\load_cnt[2]~q ),
	.datac(!\load_cnt[1]~q ),
	.datad(!\load_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\load_cnt[6]~q ),
	.datab(!\load_cnt[5]~q ),
	.datac(!\load_cnt[4]~q ),
	.datad(!\LessThan1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~1 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt[6]~1 (
	.dataa(!clk_ena),
	.datab(!dreg_11),
	.datac(!always91),
	.datad(!always9),
	.datae(!tx_rden_mii),
	.dataf(!\LessThan1~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt[6]~1 .extended_lut = "off";
defparam \load_cnt[6]~1 .lut_mask = 64'hDFFFFFFF1FFFFFFF;
defparam \load_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt[6]~2 (
	.dataa(!Selector4),
	.datab(!\Selector4~3_combout ),
	.datac(!\Selector1~4_combout ),
	.datad(!\Selector0~7_combout ),
	.datae(!\Selector0~5_combout ),
	.dataf(!\load_cnt[6]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt[6]~2 .extended_lut = "off";
defparam \load_cnt[6]~2 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \load_cnt[6]~2 .shared_arith = "off";

dffeas \load_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[0]~q ),
	.prn(vcc));
defparam \load_cnt[0] .is_wysiwyg = "true";
defparam \load_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h00000000000000FF;
defparam \Add3~21 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt~7 (
	.dataa(!\load_cnt_reg[1]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~21_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~7 .extended_lut = "off";
defparam \load_cnt~7 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~7 .shared_arith = "off";

dffeas \load_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[1]~q ),
	.prn(vcc));
defparam \load_cnt[1] .is_wysiwyg = "true";
defparam \load_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt~6 (
	.dataa(!\load_cnt_reg[2]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~17_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~6 .extended_lut = "off";
defparam \load_cnt~6 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~6 .shared_arith = "off";

dffeas \load_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[2]~q ),
	.prn(vcc));
defparam \load_cnt[2] .is_wysiwyg = "true";
defparam \load_cnt[2] .power_up = "low";

cyclonev_lcell_comb \load_cnt~5 (
	.dataa(!\load_cnt_reg[3]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~5 .extended_lut = "off";
defparam \load_cnt~5 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~5 .shared_arith = "off";

dffeas \load_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[3]~q ),
	.prn(vcc));
defparam \load_cnt[3] .is_wysiwyg = "true";
defparam \load_cnt[3] .power_up = "low";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\load_cnt[6]~q ),
	.datab(!\load_cnt[3]~q ),
	.datac(!\load_cnt[2]~q ),
	.datad(!\load_cnt[5]~q ),
	.datae(!\load_cnt[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!eop_sft_0),
	.datab(!col_int),
	.datac(!\state.STM_TYP_WAIT_END~q ),
	.datad(!\state.STM_TYP_COPY~q ),
	.datae(!\LessThan0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \Selector2~0 .shared_arith = "off";

dffeas \state.STM_TYP_WAIT_END (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_WAIT_END~q ),
	.prn(vcc));
defparam \state.STM_TYP_WAIT_END .is_wysiwyg = "true";
defparam \state.STM_TYP_WAIT_END .power_up = "low";

cyclonev_lcell_comb \Selector7~5 (
	.dataa(!eop_sft_0),
	.datab(!col_int),
	.datac(!\state.STM_TYP_WAIT_END~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~5 .extended_lut = "off";
defparam \Selector7~5 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Selector7~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~1_sumout ),
	.cout(\Add2~2 ),
	.shareout());
defparam \Add2~1 .extended_lut = "off";
defparam \Add2~1 .lut_mask = 64'h00000000000000FF;
defparam \Add2~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~0 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~1_sumout ),
	.datae(!\Add2~1_sumout ),
	.dataf(!\Add0~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~0 .extended_lut = "off";
defparam \wait_col_cnt~0 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \wait_col_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!transmit_cnt_0),
	.datab(!transmit_cnt_1),
	.datac(!transmit_cnt_2),
	.datad(!\load_cnt_reg[0]~q ),
	.datae(!\load_cnt_reg[1]~q ),
	.dataf(!\load_cnt_reg[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'h6996966996696996;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~2 (
	.dataa(!transmit_cnt_3),
	.datab(!transmit_cnt_4),
	.datac(!transmit_cnt_5),
	.datad(!\load_cnt_reg[3]~q ),
	.datae(!\load_cnt_reg[4]~q ),
	.dataf(!\load_cnt_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~2 .extended_lut = "off";
defparam \Equal1~2 .lut_mask = 64'h6996966996696996;
defparam \Equal1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~2 (
	.dataa(!eop_sft_0),
	.datab(!col_int),
	.datac(!\state.STM_TYP_COPY~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~2 .extended_lut = "off";
defparam \Selector1~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Selector1~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector1~3 (
	.dataa(!\state.STM_TYP_RETRANSMIT~q ),
	.datab(!\Equal1~0_combout ),
	.datac(!\Equal1~1_combout ),
	.datad(!\Equal1~2_combout ),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\Selector1~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~3 .extended_lut = "off";
defparam \Selector1~3 .lut_mask = 64'hFFFFDFFFFFFFFFFF;
defparam \Selector1~3 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add2~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~25_sumout ),
	.cout(\Add2~26 ),
	.shareout());
defparam \Add2~25 .extended_lut = "off";
defparam \Add2~25 .lut_mask = 64'h00000000000000FF;
defparam \Add2~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~8 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~25_sumout ),
	.datae(!\Add2~25_sumout ),
	.dataf(!\Add0~25_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~8 .extended_lut = "off";
defparam \wait_col_cnt~8 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \wait_col_cnt~8 .shared_arith = "off";

dffeas \wait_col_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~8_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[1]~q ),
	.prn(vcc));
defparam \wait_col_cnt[1] .is_wysiwyg = "true";
defparam \wait_col_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add2~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~21_sumout ),
	.cout(\Add2~22 ),
	.shareout());
defparam \Add2~21 .extended_lut = "off";
defparam \Add2~21 .lut_mask = 64'h00000000000000FF;
defparam \Add2~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000000000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~7 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~21_sumout ),
	.datae(!\Add2~21_sumout ),
	.dataf(!\Add0~21_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~7 .extended_lut = "off";
defparam \wait_col_cnt~7 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \wait_col_cnt~7 .shared_arith = "off";

dffeas \wait_col_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[2]~q ),
	.prn(vcc));
defparam \wait_col_cnt[2] .is_wysiwyg = "true";
defparam \wait_col_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add2~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~17_sumout ),
	.cout(\Add2~18 ),
	.shareout());
defparam \Add2~17 .extended_lut = "off";
defparam \Add2~17 .lut_mask = 64'h00000000000000FF;
defparam \Add2~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~6 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~17_sumout ),
	.datae(!\Add2~17_sumout ),
	.dataf(!\Add0~17_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~6 .extended_lut = "off";
defparam \wait_col_cnt~6 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \wait_col_cnt~6 .shared_arith = "off";

dffeas \wait_col_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[3]~q ),
	.prn(vcc));
defparam \wait_col_cnt[3] .is_wysiwyg = "true";
defparam \wait_col_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Add2~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~13_sumout ),
	.cout(\Add2~14 ),
	.shareout());
defparam \Add2~13 .extended_lut = "off";
defparam \Add2~13 .lut_mask = 64'h00000000000000FF;
defparam \Add2~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000000000FF00;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~5 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~13_sumout ),
	.datae(!\Add2~13_sumout ),
	.dataf(!\Add0~13_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~5 .extended_lut = "off";
defparam \wait_col_cnt~5 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \wait_col_cnt~5 .shared_arith = "off";

dffeas \wait_col_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[4]~q ),
	.prn(vcc));
defparam \wait_col_cnt[4] .is_wysiwyg = "true";
defparam \wait_col_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Add2~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~9_sumout ),
	.cout(\Add2~10 ),
	.shareout());
defparam \Add2~9 .extended_lut = "off";
defparam \Add2~9 .lut_mask = 64'h00000000000000FF;
defparam \Add2~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~4 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~9_sumout ),
	.datae(!\Add2~9_sumout ),
	.dataf(!\Add0~9_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~4 .extended_lut = "off";
defparam \wait_col_cnt~4 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \wait_col_cnt~4 .shared_arith = "off";

dffeas \wait_col_cnt[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[5]~q ),
	.prn(vcc));
defparam \wait_col_cnt[5] .is_wysiwyg = "true";
defparam \wait_col_cnt[5] .power_up = "low";

cyclonev_lcell_comb \Add2~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\wait_col_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add2~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add2~5_sumout ),
	.cout(),
	.shareout());
defparam \Add2~5 .extended_lut = "off";
defparam \Add2~5 .lut_mask = 64'h00000000000000FF;
defparam \Add2~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt~3 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\Selector1~4_combout ),
	.datac(!\Selector7~5_combout ),
	.datad(!\Add1~5_sumout ),
	.datae(!\Add2~5_sumout ),
	.dataf(!\Add0~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt~3 .extended_lut = "off";
defparam \wait_col_cnt~3 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \wait_col_cnt~3 .shared_arith = "off";

dffeas \wait_col_cnt[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[6]~q ),
	.prn(vcc));
defparam \wait_col_cnt[6] .is_wysiwyg = "true";
defparam \wait_col_cnt[6] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\wait_col_cnt[6]~q ),
	.datab(!\wait_col_cnt[5]~q ),
	.datac(!\wait_col_cnt[4]~q ),
	.datad(!\wait_col_cnt[3]~q ),
	.datae(!\wait_col_cnt[2]~q ),
	.dataf(!\wait_col_cnt[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~6 (
	.dataa(!eop_sft_0),
	.datab(!\state.STM_TYP_COPY~q ),
	.datac(!\state.STM_TYP_WAIT_COL~q ),
	.datad(!\wait_col_cnt[0]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~6 .extended_lut = "off";
defparam \Selector7~6 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Selector7~6 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt[6]~1 (
	.dataa(!clk_ena),
	.datab(!stateSTM_TYP_WAIT_COL_1),
	.datac(!col_int),
	.datad(!\Selector7~6_combout ),
	.datae(!\Selector7~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt[6]~1 .extended_lut = "off";
defparam \wait_col_cnt[6]~1 .lut_mask = 64'hFFFFEFFFFFFFEFFF;
defparam \wait_col_cnt[6]~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_col_cnt[6]~2 (
	.dataa(!stateSTM_TYP_WAIT_COL_1),
	.datab(!\col_reg~q ),
	.datac(!Selector1),
	.datad(!\Selector1~3_combout ),
	.datae(!\wait_col_cnt[6]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_col_cnt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_col_cnt[6]~2 .extended_lut = "off";
defparam \wait_col_cnt[6]~2 .lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam \wait_col_cnt[6]~2 .shared_arith = "off";

dffeas \wait_col_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_col_cnt~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wait_col_cnt[6]~2_combout ),
	.q(\wait_col_cnt[0]~q ),
	.prn(vcc));
defparam \wait_col_cnt[0] .is_wysiwyg = "true";
defparam \wait_col_cnt[0] .power_up = "low";

cyclonev_lcell_comb \always0~4 (
	.dataa(!eop_sft_0),
	.datab(!\state.STM_TYP_COPY~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~4 .extended_lut = "off";
defparam \always0~4 .lut_mask = 64'h7777777777777777;
defparam \always0~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~3 (
	.dataa(!clk_ena),
	.datab(!eop_sft_0),
	.datac(!stateSTM_TYP_WAIT_COL_1),
	.datad(!col_int),
	.datae(!\state.STM_TYP_WAIT_END~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~3 .extended_lut = "off";
defparam \Selector7~3 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \Selector7~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector7~4 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\wait_col_cnt[0]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(!\always0~4_combout ),
	.dataf(!\Selector7~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector7~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector7~4 .extended_lut = "off";
defparam \Selector7~4 .lut_mask = 64'hFFBFFFFFFFFFFFFF;
defparam \Selector7~4 .shared_arith = "off";

dffeas \state.STM_TYP_WAIT_COL (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector7~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_WAIT_COL~q ),
	.prn(vcc));
defparam \state.STM_TYP_WAIT_COL .is_wysiwyg = "true";
defparam \state.STM_TYP_WAIT_COL .power_up = "low";

cyclonev_lcell_comb \Add6~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~13_sumout ),
	.cout(\Add6~14 ),
	.shareout());
defparam \Add6~13 .extended_lut = "off";
defparam \Add6~13 .lut_mask = 64'h00000000000000FF;
defparam \Add6~13 .shared_arith = "off";

cyclonev_lcell_comb \always14~0 (
	.dataa(!clk_ena),
	.datab(!\state.STM_TYP_BACK_OFF~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always14~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always14~0 .extended_lut = "off";
defparam \always14~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \always14~0 .shared_arith = "off";

cyclonev_lcell_comb \Add6~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~1_sumout ),
	.cout(\Add6~2 ),
	.shareout());
defparam \Add6~1 .extended_lut = "off";
defparam \Add6~1 .lut_mask = 64'h00000000000000FF;
defparam \Add6~1 .shared_arith = "off";

cyclonev_lcell_comb \Add6~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~61_sumout ),
	.cout(\Add6~62 ),
	.shareout());
defparam \Add6~61 .extended_lut = "off";
defparam \Add6~61 .lut_mask = 64'h00000000000000FF;
defparam \Add6~61 .shared_arith = "off";

dffeas \back_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~61_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[4]~q ),
	.prn(vcc));
defparam \back_cnt[4] .is_wysiwyg = "true";
defparam \back_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Add6~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~57_sumout ),
	.cout(\Add6~58 ),
	.shareout());
defparam \Add6~57 .extended_lut = "off";
defparam \Add6~57 .lut_mask = 64'h00000000000000FF;
defparam \Add6~57 .shared_arith = "off";

dffeas \back_cnt[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~57_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[5]~q ),
	.prn(vcc));
defparam \back_cnt[5] .is_wysiwyg = "true";
defparam \back_cnt[5] .power_up = "low";

cyclonev_lcell_comb \Add6~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~53_sumout ),
	.cout(\Add6~54 ),
	.shareout());
defparam \Add6~53 .extended_lut = "off";
defparam \Add6~53 .lut_mask = 64'h00000000000000FF;
defparam \Add6~53 .shared_arith = "off";

dffeas \back_cnt[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~53_sumout ),
	.asdata(\U_LFSR|z_reg[0]~q ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[6]~q ),
	.prn(vcc));
defparam \back_cnt[6] .is_wysiwyg = "true";
defparam \back_cnt[6] .power_up = "low";

cyclonev_lcell_comb \Add6~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~49_sumout ),
	.cout(\Add6~50 ),
	.shareout());
defparam \Add6~49 .extended_lut = "off";
defparam \Add6~49 .lut_mask = 64'h00000000000000FF;
defparam \Add6~49 .shared_arith = "off";

cyclonev_lcell_comb \wait_late~0 (
	.dataa(!dreg_1),
	.datab(!col_int),
	.datac(!\state.STM_TYP_WAIT_COL~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_late~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_late~0 .extended_lut = "off";
defparam \wait_late~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \wait_late~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_late~1 (
	.dataa(!\state.STM_TYP_WAIT_COL~q ),
	.datab(!\wait_col_cnt[0]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!crs),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_late~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_late~1 .extended_lut = "off";
defparam \wait_late~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \wait_late~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_late~2 (
	.dataa(!eop_sft_0),
	.datab(!col_int),
	.datac(!\state.STM_TYP_WAIT_END~q ),
	.datad(!\state.STM_TYP_COPY~q ),
	.datae(!\LessThan0~0_combout ),
	.dataf(!\wait_late~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_late~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_late~2 .extended_lut = "off";
defparam \wait_late~2 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \wait_late~2 .shared_arith = "off";

cyclonev_lcell_comb \wait_late~3 (
	.dataa(!\state.STM_TYP_IDLE~q ),
	.datab(!\Selector0~2_combout ),
	.datac(!\wait_late~q ),
	.datad(!crs),
	.datae(!\wait_late~0_combout ),
	.dataf(!\wait_late~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_late~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_late~3 .extended_lut = "off";
defparam \wait_late~3 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \wait_late~3 .shared_arith = "off";

dffeas wait_late(
	.clk(mac_tx_clock_connection_clk),
	.d(\wait_late~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_late~q ),
	.prn(vcc));
defparam wait_late.is_wysiwyg = "true";
defparam wait_late.power_up = "low";

cyclonev_lcell_comb \Selector6~2 (
	.dataa(!\state.STM_TYP_WAIT_COL~q ),
	.datab(!\wait_col_cnt[0]~q ),
	.datac(!\wait_late~q ),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~2 .extended_lut = "off";
defparam \Selector6~2 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \Selector6~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~8 (
	.dataa(!\state.STM_TYP_RETRANSMIT~q ),
	.datab(!\Equal1~1_combout ),
	.datac(!\Equal1~2_combout ),
	.datad(!\state.STM_TYP_COPY~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~8 .extended_lut = "off";
defparam \Selector6~8 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \Selector6~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~6 (
	.dataa(!\state.STM_TYP_RETRANSMIT~q ),
	.datab(!\Equal1~0_combout ),
	.datac(!\Selector6~2_combout ),
	.datad(!q_b_9),
	.datae(!stateSTM_TYP_RETRANSMIT_SHORT),
	.dataf(!\Selector6~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~6 .extended_lut = "off";
defparam \Selector6~6 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Selector6~6 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt~0 (
	.dataa(!stateSTM_TYP_RETRANSMIT_SHORT),
	.datab(!\state.STM_TYP_RETRANSMIT~q ),
	.datac(!\state.STM_TYP_COPY~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt~0 .extended_lut = "off";
defparam \retrans_cnt~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \retrans_cnt~0 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt~7 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~6_combout ),
	.datae(!\retrans_cnt[0]~q ),
	.dataf(!\retrans_cnt~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt~7 .extended_lut = "off";
defparam \retrans_cnt~7 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \retrans_cnt~7 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt[3]~2 (
	.dataa(!\col_reg~q ),
	.datab(!\state.STM_TYP_IDLE~q ),
	.datac(!\state.STM_TYP_FLUSH~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt[3]~2 .extended_lut = "off";
defparam \retrans_cnt[3]~2 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \retrans_cnt[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt[3]~3 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~6_combout ),
	.datae(!\retrans_cnt~0_combout ),
	.dataf(!\retrans_cnt[3]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt[3]~3 .extended_lut = "off";
defparam \retrans_cnt[3]~3 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \retrans_cnt[3]~3 .shared_arith = "off";

dffeas \retrans_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\retrans_cnt~7_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\retrans_cnt[3]~3_combout ),
	.q(\retrans_cnt[0]~q ),
	.prn(vcc));
defparam \retrans_cnt[0] .is_wysiwyg = "true";
defparam \retrans_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add5~3 (
	.dataa(!\retrans_cnt[1]~q ),
	.datab(!\retrans_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~3 .extended_lut = "off";
defparam \Add5~3 .lut_mask = 64'h6666666666666666;
defparam \Add5~3 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt~6 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~6_combout ),
	.datae(!\retrans_cnt~0_combout ),
	.dataf(!\Add5~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt~6 .extended_lut = "off";
defparam \retrans_cnt~6 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \retrans_cnt~6 .shared_arith = "off";

dffeas \retrans_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\retrans_cnt~6_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\retrans_cnt[3]~3_combout ),
	.q(\retrans_cnt[1]~q ),
	.prn(vcc));
defparam \retrans_cnt[1] .is_wysiwyg = "true";
defparam \retrans_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add5~2 (
	.dataa(!\retrans_cnt[2]~q ),
	.datab(!\retrans_cnt[1]~q ),
	.datac(!\retrans_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~2 .extended_lut = "off";
defparam \Add5~2 .lut_mask = 64'h9696969696969696;
defparam \Add5~2 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt~5 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~6_combout ),
	.datae(!\retrans_cnt~0_combout ),
	.dataf(!\Add5~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt~5 .extended_lut = "off";
defparam \retrans_cnt~5 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \retrans_cnt~5 .shared_arith = "off";

dffeas \retrans_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\retrans_cnt~5_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\retrans_cnt[3]~3_combout ),
	.q(\retrans_cnt[2]~q ),
	.prn(vcc));
defparam \retrans_cnt[2] .is_wysiwyg = "true";
defparam \retrans_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add5~1 (
	.dataa(!\retrans_cnt[3]~q ),
	.datab(!\retrans_cnt[2]~q ),
	.datac(!\retrans_cnt[1]~q ),
	.datad(!\retrans_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~1 .extended_lut = "off";
defparam \Add5~1 .lut_mask = 64'h6996699669966996;
defparam \Add5~1 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt~4 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~6_combout ),
	.datae(!\retrans_cnt~0_combout ),
	.dataf(!\Add5~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt~4 .extended_lut = "off";
defparam \retrans_cnt~4 .lut_mask = 64'hFFFFFF7FFFFFFFFF;
defparam \retrans_cnt~4 .shared_arith = "off";

dffeas \retrans_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\retrans_cnt~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\retrans_cnt[3]~3_combout ),
	.q(\retrans_cnt[3]~q ),
	.prn(vcc));
defparam \retrans_cnt[3] .is_wysiwyg = "true";
defparam \retrans_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Equal3~0 (
	.dataa(!\retrans_cnt[2]~q ),
	.datab(!\retrans_cnt[1]~q ),
	.datac(!\retrans_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal3~0 .extended_lut = "off";
defparam \Equal3~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~9 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\Equal3~0_combout ),
	.datad(!\U_LFSR|z_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~9 .extended_lut = "off";
defparam \back_cnt~9 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \back_cnt~9 .shared_arith = "off";

dffeas \back_cnt[7] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~49_sumout ),
	.asdata(\back_cnt~9_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[7]~q ),
	.prn(vcc));
defparam \back_cnt[7] .is_wysiwyg = "true";
defparam \back_cnt[7] .power_up = "low";

cyclonev_lcell_comb \Add6~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~45_sumout ),
	.cout(\Add6~46 ),
	.shareout());
defparam \Add6~45 .extended_lut = "off";
defparam \Add6~45 .lut_mask = 64'h00000000000000FF;
defparam \Add6~45 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~8 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\retrans_cnt[1]~q ),
	.datae(!\U_LFSR|z_reg[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~8 .extended_lut = "off";
defparam \back_cnt~8 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \back_cnt~8 .shared_arith = "off";

dffeas \back_cnt[8] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~45_sumout ),
	.asdata(\back_cnt~8_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[8]~q ),
	.prn(vcc));
defparam \back_cnt[8] .is_wysiwyg = "true";
defparam \back_cnt[8] .power_up = "low";

cyclonev_lcell_comb \Add6~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~41_sumout ),
	.cout(\Add6~42 ),
	.shareout());
defparam \Add6~41 .extended_lut = "off";
defparam \Add6~41 .lut_mask = 64'h00000000000000FF;
defparam \Add6~41 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~7 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\retrans_cnt[1]~q ),
	.datae(!\retrans_cnt[0]~q ),
	.dataf(!\U_LFSR|z_reg[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~7 .extended_lut = "off";
defparam \back_cnt~7 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \back_cnt~7 .shared_arith = "off";

dffeas \back_cnt[9] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~41_sumout ),
	.asdata(\back_cnt~7_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[9]~q ),
	.prn(vcc));
defparam \back_cnt[9] .is_wysiwyg = "true";
defparam \back_cnt[9] .power_up = "low";

cyclonev_lcell_comb \Add6~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~37_sumout ),
	.cout(\Add6~38 ),
	.shareout());
defparam \Add6~37 .extended_lut = "off";
defparam \Add6~37 .lut_mask = 64'h00000000000000FF;
defparam \Add6~37 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~6 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\U_LFSR|z_reg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~6 .extended_lut = "off";
defparam \back_cnt~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \back_cnt~6 .shared_arith = "off";

dffeas \back_cnt[10] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~37_sumout ),
	.asdata(\back_cnt~6_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[10]~q ),
	.prn(vcc));
defparam \back_cnt[10] .is_wysiwyg = "true";
defparam \back_cnt[10] .power_up = "low";

cyclonev_lcell_comb \Add6~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~33_sumout ),
	.cout(\Add6~34 ),
	.shareout());
defparam \Add6~33 .extended_lut = "off";
defparam \Add6~33 .lut_mask = 64'h00000000000000FF;
defparam \Add6~33 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~5 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\retrans_cnt[1]~q ),
	.datae(!\retrans_cnt[0]~q ),
	.dataf(!\U_LFSR|z_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~5 .extended_lut = "off";
defparam \back_cnt~5 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \back_cnt~5 .shared_arith = "off";

dffeas \back_cnt[11] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~33_sumout ),
	.asdata(\back_cnt~5_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[11]~q ),
	.prn(vcc));
defparam \back_cnt[11] .is_wysiwyg = "true";
defparam \back_cnt[11] .power_up = "low";

cyclonev_lcell_comb \Add6~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~29_sumout ),
	.cout(\Add6~30 ),
	.shareout());
defparam \Add6~29 .extended_lut = "off";
defparam \Add6~29 .lut_mask = 64'h00000000000000FF;
defparam \Add6~29 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~4 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\retrans_cnt[1]~q ),
	.datae(!\U_LFSR|z_reg[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~4 .extended_lut = "off";
defparam \back_cnt~4 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \back_cnt~4 .shared_arith = "off";

dffeas \back_cnt[12] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~29_sumout ),
	.asdata(\back_cnt~4_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[12]~q ),
	.prn(vcc));
defparam \back_cnt[12] .is_wysiwyg = "true";
defparam \back_cnt[12] .power_up = "low";

cyclonev_lcell_comb \Add6~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~25_sumout ),
	.cout(\Add6~26 ),
	.shareout());
defparam \Add6~25 .extended_lut = "off";
defparam \Add6~25 .lut_mask = 64'h00000000000000FF;
defparam \Add6~25 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~3 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\retrans_cnt[1]~q ),
	.datae(!\retrans_cnt[0]~q ),
	.dataf(!\U_LFSR|z_reg[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~3 .extended_lut = "off";
defparam \back_cnt~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \back_cnt~3 .shared_arith = "off";

dffeas \back_cnt[13] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~25_sumout ),
	.asdata(\back_cnt~3_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[13]~q ),
	.prn(vcc));
defparam \back_cnt[13] .is_wysiwyg = "true";
defparam \back_cnt[13] .power_up = "low";

cyclonev_lcell_comb \Add6~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~21_sumout ),
	.cout(\Add6~22 ),
	.shareout());
defparam \Add6~21 .extended_lut = "off";
defparam \Add6~21 .lut_mask = 64'h00000000000000FF;
defparam \Add6~21 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~2 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(gnd),
	.datad(!\U_LFSR|z_reg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~2 .extended_lut = "off";
defparam \back_cnt~2 .lut_mask = 64'h77FF77FF77FF77FF;
defparam \back_cnt~2 .shared_arith = "off";

dffeas \back_cnt[14] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~21_sumout ),
	.asdata(\back_cnt~2_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[14]~q ),
	.prn(vcc));
defparam \back_cnt[14] .is_wysiwyg = "true";
defparam \back_cnt[14] .power_up = "low";

cyclonev_lcell_comb \Add6~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~17_sumout ),
	.cout(),
	.shareout());
defparam \Add6~17 .extended_lut = "off";
defparam \Add6~17 .lut_mask = 64'h00000000000000FF;
defparam \Add6~17 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~1 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(gnd),
	.datad(!\Equal3~0_combout ),
	.datae(!\U_LFSR|z_reg[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~1 .extended_lut = "off";
defparam \back_cnt~1 .lut_mask = 64'hFF77FFFFFF77FFFF;
defparam \back_cnt~1 .shared_arith = "off";

dffeas \back_cnt[15] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~17_sumout ),
	.asdata(\back_cnt~1_combout ),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[15]~q ),
	.prn(vcc));
defparam \back_cnt[15] .is_wysiwyg = "true";
defparam \back_cnt[15] .power_up = "low";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!\back_cnt[15]~q ),
	.datab(!\back_cnt[14]~q ),
	.datac(!\back_cnt[13]~q ),
	.datad(!\back_cnt[12]~q ),
	.datae(!\back_cnt[11]~q ),
	.dataf(!\back_cnt[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~2 (
	.dataa(!\back_cnt[9]~q ),
	.datab(!\back_cnt[8]~q ),
	.datac(!\back_cnt[7]~q ),
	.datad(!\back_cnt[6]~q ),
	.datae(!\back_cnt[5]~q ),
	.dataf(!\back_cnt[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~2 .extended_lut = "off";
defparam \Equal2~2 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal2~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~3 (
	.dataa(!\Equal2~0_combout ),
	.datab(!\Equal2~1_combout ),
	.datac(!\Equal2~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~3 .extended_lut = "off";
defparam \Equal2~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal2~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~7 (
	.dataa(!\state.STM_TYP_RETRANSMIT~q ),
	.datab(!\Equal1~2_combout ),
	.datac(!\state.STM_TYP_COPY~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~7 .extended_lut = "off";
defparam \Selector6~7 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Selector6~7 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~5 (
	.dataa(!\state.STM_TYP_RETRANSMIT~q ),
	.datab(!\Equal1~0_combout ),
	.datac(!\Equal1~1_combout ),
	.datad(!q_b_9),
	.datae(!stateSTM_TYP_RETRANSMIT_SHORT),
	.dataf(!\Selector6~7_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~5 .extended_lut = "off";
defparam \Selector6~5 .lut_mask = 64'hFFFFEFFFFFFFFFFF;
defparam \Selector6~5 .shared_arith = "off";

cyclonev_lcell_comb \back_cnt~0 (
	.dataa(!clk_ena),
	.datab(!col_int),
	.datac(!\state.STM_TYP_BACK_OFF~q ),
	.datad(!\Equal2~3_combout ),
	.datae(!\Selector6~2_combout ),
	.dataf(!\Selector6~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\back_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \back_cnt~0 .extended_lut = "off";
defparam \back_cnt~0 .lut_mask = 64'hFF7FFFFFF777FFFF;
defparam \back_cnt~0 .shared_arith = "off";

dffeas \back_cnt[0] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~13_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[0]~q ),
	.prn(vcc));
defparam \back_cnt[0] .is_wysiwyg = "true";
defparam \back_cnt[0] .power_up = "low";

cyclonev_lcell_comb \Add6~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~9_sumout ),
	.cout(\Add6~10 ),
	.shareout());
defparam \Add6~9 .extended_lut = "off";
defparam \Add6~9 .lut_mask = 64'h00000000000000FF;
defparam \Add6~9 .shared_arith = "off";

dffeas \back_cnt[1] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~9_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[1]~q ),
	.prn(vcc));
defparam \back_cnt[1] .is_wysiwyg = "true";
defparam \back_cnt[1] .power_up = "low";

cyclonev_lcell_comb \Add6~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\back_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add6~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add6~5_sumout ),
	.cout(\Add6~6 ),
	.shareout());
defparam \Add6~5 .extended_lut = "off";
defparam \Add6~5 .lut_mask = 64'h00000000000000FF;
defparam \Add6~5 .shared_arith = "off";

dffeas \back_cnt[2] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~5_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[2]~q ),
	.prn(vcc));
defparam \back_cnt[2] .is_wysiwyg = "true";
defparam \back_cnt[2] .power_up = "low";

dffeas \back_cnt[3] (
	.clk(mac_tx_clock_connection_clk),
	.d(\Add6~1_sumout ),
	.asdata(GND_port),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always14~0_combout ),
	.ena(\back_cnt~0_combout ),
	.q(\back_cnt[3]~q ),
	.prn(vcc));
defparam \back_cnt[3] .is_wysiwyg = "true";
defparam \back_cnt[3] .power_up = "low";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\back_cnt[3]~q ),
	.datab(!\back_cnt[2]~q ),
	.datac(!\back_cnt[1]~q ),
	.datad(!\back_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~1 (
	.dataa(!\state.STM_TYP_BACK_OFF~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\Equal2~1_combout ),
	.datad(!\Equal2~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~1 .extended_lut = "off";
defparam \Selector6~1 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Selector6~1 .shared_arith = "off";

cyclonev_lcell_comb \Add5~0 (
	.dataa(!\retrans_cnt[4]~q ),
	.datab(!\retrans_cnt[3]~q ),
	.datac(!\retrans_cnt[2]~q ),
	.datad(!\retrans_cnt[1]~q ),
	.datae(!\retrans_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add5~0 .extended_lut = "off";
defparam \Add5~0 .lut_mask = 64'h9669699696696996;
defparam \Add5~0 .shared_arith = "off";

cyclonev_lcell_comb \retrans_cnt~1 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~6_combout ),
	.datae(!\Add5~0_combout ),
	.dataf(!\retrans_cnt~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\retrans_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \retrans_cnt~1 .extended_lut = "off";
defparam \retrans_cnt~1 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \retrans_cnt~1 .shared_arith = "off";

dffeas \retrans_cnt[4] (
	.clk(mac_tx_clock_connection_clk),
	.d(\retrans_cnt~1_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\retrans_cnt[3]~3_combout ),
	.q(\retrans_cnt[4]~q ),
	.prn(vcc));
defparam \retrans_cnt[4] .is_wysiwyg = "true";
defparam \retrans_cnt[4] .power_up = "low";

cyclonev_lcell_comb \always16~0 (
	.dataa(!\state.STM_TYP_FLUSH~q ),
	.datab(!\retrans_cnt[4]~q ),
	.datac(!\retrans_cnt[3]~q ),
	.datad(!\Equal3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always16~0 .extended_lut = "off";
defparam \always16~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \always16~0 .shared_arith = "off";

dffeas excess_col_int(
	.clk(mac_tx_clock_connection_clk),
	.d(\always16~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\excess_col_int~q ),
	.prn(vcc));
defparam excess_col_int.is_wysiwyg = "true";
defparam excess_col_int.power_up = "low";

cyclonev_lcell_comb \Selector0~2 (
	.dataa(!clk_ena),
	.datab(!dreg_11),
	.datac(!always91),
	.datad(!always9),
	.datae(!\excess_col_int~q ),
	.dataf(!tx_rden_mii),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~2 .extended_lut = "off";
defparam \Selector0~2 .lut_mask = 64'hFFFFFFFFFFFFFFB8;
defparam \Selector0~2 .shared_arith = "off";

cyclonev_lcell_comb \col_reg~0 (
	.dataa(!\col_reg~q ),
	.datab(!\state.STM_TYP_IDLE~q ),
	.datac(!\Selector0~2_combout ),
	.datad(!\wait_late~q ),
	.datae(!\Selector0~5_combout ),
	.dataf(!\Selector6~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\col_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \col_reg~0 .extended_lut = "off";
defparam \col_reg~0 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \col_reg~0 .shared_arith = "off";

dffeas col_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(\col_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\col_reg~q ),
	.prn(vcc));
defparam col_reg.is_wysiwyg = "true";
defparam col_reg.power_up = "low";

cyclonev_lcell_comb \Selector1~4 (
	.dataa(!dreg_11),
	.datab(!\col_reg~q ),
	.datac(!always92),
	.datad(!tx_rden_mii),
	.datae(!\Selector1~0_combout ),
	.dataf(!\Selector1~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector1~4 .extended_lut = "off";
defparam \Selector1~4 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \Selector1~4 .shared_arith = "off";

dffeas \state.STM_TYP_COPY (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector1~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_COPY~q ),
	.prn(vcc));
defparam \state.STM_TYP_COPY .is_wysiwyg = "true";
defparam \state.STM_TYP_COPY .power_up = "low";

cyclonev_lcell_comb \load_cnt_reg~0 (
	.dataa(!eop_sft_0),
	.datab(!col_int),
	.datac(!\state.STM_TYP_COPY~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt_reg~0 .extended_lut = "off";
defparam \load_cnt_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \load_cnt_reg~0 .shared_arith = "off";

dffeas \load_cnt_reg[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[5]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[5]~q ),
	.prn(vcc));
defparam \load_cnt_reg[5] .is_wysiwyg = "true";
defparam \load_cnt_reg[5] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt~3 (
	.dataa(!\load_cnt_reg[5]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~5_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~3 .extended_lut = "off";
defparam \load_cnt~3 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~3 .shared_arith = "off";

dffeas \load_cnt[5] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~3_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[5]~q ),
	.prn(vcc));
defparam \load_cnt[5] .is_wysiwyg = "true";
defparam \load_cnt[5] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\load_cnt[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \load_cnt~0 (
	.dataa(!\load_cnt_reg[6]~q ),
	.datab(!Selector4),
	.datac(!short_frm1),
	.datad(!Selector1),
	.datae(!Selector5),
	.dataf(!\Add3~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\load_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \load_cnt~0 .extended_lut = "off";
defparam \load_cnt~0 .lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam \load_cnt~0 .shared_arith = "off";

dffeas \load_cnt[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(\Selector0~6_combout ),
	.sload(gnd),
	.ena(\load_cnt[6]~2_combout ),
	.q(\load_cnt[6]~q ),
	.prn(vcc));
defparam \load_cnt[6] .is_wysiwyg = "true";
defparam \load_cnt[6] .power_up = "low";

dffeas \load_cnt_reg[6] (
	.clk(mac_tx_clock_connection_clk),
	.d(\load_cnt[6]~q ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_cnt_reg~0_combout ),
	.q(\load_cnt_reg[6]~q ),
	.prn(vcc));
defparam \load_cnt_reg[6] .is_wysiwyg = "true";
defparam \load_cnt_reg[6] .power_up = "low";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!transmit_cnt_6),
	.datab(!\load_cnt_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'h6666666666666666;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector4~2 (
	.dataa(!\state.STM_TYP_RETRANSMIT~q ),
	.datab(!\Equal1~0_combout ),
	.datac(!\Equal1~1_combout ),
	.datad(!\Equal1~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector4~2 .extended_lut = "off";
defparam \Selector4~2 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \Selector4~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~3 (
	.dataa(!q_b_9),
	.datab(!stateSTM_TYP_RETRANSMIT_SHORT),
	.datac(!\state.STM_TYP_COPY~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~3 .extended_lut = "off";
defparam \Selector6~3 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Selector6~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector6~4 (
	.dataa(!col_int),
	.datab(!\Selector4~2_combout ),
	.datac(!\Selector6~1_combout ),
	.datad(!\Selector6~2_combout ),
	.datae(!\Selector6~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector6~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector6~4 .extended_lut = "off";
defparam \Selector6~4 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \Selector6~4 .shared_arith = "off";

dffeas \state.STM_TYP_BACK_OFF (
	.clk(mac_tx_clock_connection_clk),
	.d(\Selector6~4_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.STM_TYP_BACK_OFF~q ),
	.prn(vcc));
defparam \state.STM_TYP_BACK_OFF .is_wysiwyg = "true";
defparam \state.STM_TYP_BACK_OFF .power_up = "low";

cyclonev_lcell_comb \Selector0~3 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(!\wait_col_cnt[0]~q ),
	.datad(!\wait_late~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~3 .extended_lut = "off";
defparam \Selector0~3 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \Selector0~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~4 (
	.dataa(!dreg_1),
	.datab(!eop_sft_0),
	.datac(!short_frm1),
	.datad(!\state.STM_TYP_IDLE~q ),
	.datae(!\state.STM_TYP_FLUSH~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~4 .extended_lut = "off";
defparam \Selector0~4 .lut_mask = 64'hFFFFFDFFFFFFFDFF;
defparam \Selector0~4 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~5 (
	.dataa(!\state.STM_TYP_BACK_OFF~q ),
	.datab(!\Equal2~0_combout ),
	.datac(!\Equal2~1_combout ),
	.datad(!\Equal2~2_combout ),
	.datae(!\Selector0~3_combout ),
	.dataf(!\Selector0~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~5 .extended_lut = "off";
defparam \Selector0~5 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Selector0~5 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~8 (
	.dataa(!\state.STM_TYP_IDLE~q ),
	.datab(!dreg_11),
	.datac(!\excess_col_int~q ),
	.datad(!tx_rden_mii),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~8 .extended_lut = "off";
defparam \Selector0~8 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \Selector0~8 .shared_arith = "off";

cyclonev_lcell_comb \Selector0~6 (
	.dataa(!\Selector0~5_combout ),
	.datab(!clk_ena),
	.datac(!dreg_11),
	.datad(!always91),
	.datae(!always9),
	.dataf(!\Selector0~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector0~6 .extended_lut = "off";
defparam \Selector0~6 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Selector0~6 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~1 (
	.dataa(!q_b_9),
	.datab(!stateSTM_TYP_RETRANSMIT_SHORT),
	.datac(!col_int),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~1 .extended_lut = "off";
defparam \Selector5~1 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \Selector5~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~3 (
	.dataa(!short_frm1),
	.datab(!clk_ena),
	.datac(!dreg_11),
	.datad(!tx_rden_mii),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~3 .extended_lut = "off";
defparam \Selector5~3 .lut_mask = 64'h53FFFFFF53FFFFFF;
defparam \Selector5~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector5~2 (
	.dataa(!Selector5),
	.datab(!\Selector5~1_combout ),
	.datac(!dreg_11),
	.datad(!always91),
	.datae(!always9),
	.dataf(!\Selector5~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector5~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector5~2 .extended_lut = "off";
defparam \Selector5~2 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \Selector5~2 .shared_arith = "off";

dffeas clk_ena_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(clk_ena),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_ena_reg~q ),
	.prn(vcc));
defparam clk_ena_reg.is_wysiwyg = "true";
defparam clk_ena_reg.power_up = "low";

cyclonev_lcell_comb \mac_ff_rden_reg~0 (
	.dataa(!tx_rden_int),
	.datab(!\mac_ff_rden_reg~q ),
	.datac(!\clk_ena_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mac_ff_rden_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mac_ff_rden_reg~0 .extended_lut = "off";
defparam \mac_ff_rden_reg~0 .lut_mask = 64'h5353535353535353;
defparam \mac_ff_rden_reg~0 .shared_arith = "off";

dffeas mac_ff_rden_reg(
	.clk(mac_tx_clock_connection_clk),
	.d(\mac_ff_rden_reg~0_combout ),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mac_ff_rden_reg~q ),
	.prn(vcc));
defparam mac_ff_rden_reg.is_wysiwyg = "true";
defparam mac_ff_rden_reg.power_up = "low";

cyclonev_lcell_comb \transmit_cnt[6]~0 (
	.dataa(!clk_ena),
	.datab(!\Selector4~1_combout ),
	.datac(!\Selector5~2_combout ),
	.datad(!\mac_ff_rden_reg~q ),
	.datae(!\Selector0~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\transmit_cnt[6]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \transmit_cnt[6]~0 .extended_lut = "off";
defparam \transmit_cnt[6]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \transmit_cnt[6]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add4~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~5_sumout ),
	.cout(\Add4~6 ),
	.shareout());
defparam \Add4~5 .extended_lut = "off";
defparam \Add4~5 .lut_mask = 64'h00000000000000FF;
defparam \Add4~5 .shared_arith = "off";

cyclonev_lcell_comb \Add4~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~9_sumout ),
	.cout(\Add4~10 ),
	.shareout());
defparam \Add4~9 .extended_lut = "off";
defparam \Add4~9 .lut_mask = 64'h00000000000000FF;
defparam \Add4~9 .shared_arith = "off";

cyclonev_lcell_comb \Add4~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~13_sumout ),
	.cout(\Add4~14 ),
	.shareout());
defparam \Add4~13 .extended_lut = "off";
defparam \Add4~13 .lut_mask = 64'h00000000000000FF;
defparam \Add4~13 .shared_arith = "off";

cyclonev_lcell_comb \Add4~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~17_sumout ),
	.cout(\Add4~18 ),
	.shareout());
defparam \Add4~17 .extended_lut = "off";
defparam \Add4~17 .lut_mask = 64'h00000000000000FF;
defparam \Add4~17 .shared_arith = "off";

cyclonev_lcell_comb \Add4~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~21_sumout ),
	.cout(\Add4~22 ),
	.shareout());
defparam \Add4~21 .extended_lut = "off";
defparam \Add4~21 .lut_mask = 64'h00000000000000FF;
defparam \Add4~21 .shared_arith = "off";

cyclonev_lcell_comb \Add4~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!transmit_cnt_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add4~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add4~25_sumout ),
	.cout(),
	.shareout());
defparam \Add4~25 .extended_lut = "off";
defparam \Add4~25 .lut_mask = 64'h00000000000000FF;
defparam \Add4~25 .shared_arith = "off";

cyclonev_lcell_comb \always9~0 (
	.dataa(!\col_reg~q ),
	.datab(!Selector1),
	.datac(!\LessThan1~1_combout ),
	.datad(!\Selector1~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always9~0 .extended_lut = "off";
defparam \always9~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \always9~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!clk_ena),
	.datab(!q_b_9),
	.datac(!stateSTM_TYP_WAIT_COL_1),
	.datad(!stateSTM_TYP_RETRANSMIT_SHORT),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~3 (
	.dataa(!\state.STM_TYP_FLUSH~q ),
	.datab(!\state.STM_TYP_WAIT_COL~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~3 .extended_lut = "off";
defparam \always0~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \always0~3 .shared_arith = "off";

cyclonev_lcell_comb \always0~5 (
	.dataa(!col_int),
	.datab(!\always0~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~5 .extended_lut = "off";
defparam \always0~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always0~5 .shared_arith = "off";

cyclonev_lcell_comb \short_frm~0 (
	.dataa(!short_frm1),
	.datab(!\state.STM_TYP_IDLE~q ),
	.datac(!\Selector0~2_combout ),
	.datad(!\Selector0~5_combout ),
	.datae(!\always0~3_combout ),
	.dataf(!\always0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\short_frm~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \short_frm~0 .extended_lut = "off";
defparam \short_frm~0 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \short_frm~0 .shared_arith = "off";

cyclonev_lcell_comb \always10~1 (
	.dataa(!Selector5),
	.datab(!clk_ena),
	.datac(!dreg_11),
	.datad(!tx_rden_mii),
	.datae(!\Selector1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~1 .extended_lut = "off";
defparam \always10~1 .lut_mask = 64'h53FFFFFF53FFFFFF;
defparam \always10~1 .shared_arith = "off";

cyclonev_lcell_comb \always10~2 (
	.dataa(!dreg_11),
	.datab(!always9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always10~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always10~2 .extended_lut = "off";
defparam \always10~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always10~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector3~1 (
	.dataa(!col_int),
	.datab(!\state.STM_TYP_WAIT_END~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector3~1 .extended_lut = "off";
defparam \Selector3~1 .lut_mask = 64'h7777777777777777;
defparam \Selector3~1 .shared_arith = "off";

dffeas crs_d(
	.clk(mac_tx_clock_connection_clk),
	.d(crs),
	.asdata(vcc),
	.clrn(altera_tse_reset_synchronizer_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clk_ena),
	.q(\crs_d~q ),
	.prn(vcc));
defparam crs_d.is_wysiwyg = "true";
defparam crs_d.power_up = "low";

cyclonev_lcell_comb \mac_ena~0 (
	.dataa(!crs),
	.datab(!\crs_d~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mac_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mac_ena~0 .extended_lut = "off";
defparam \mac_ena~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \mac_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \mac_ena~1 (
	.dataa(!\state.STM_TYP_FLUSH~q ),
	.datab(!\state.STM_TYP_BACK_OFF~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mac_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mac_ena~1 .extended_lut = "off";
defparam \mac_ena~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \mac_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \mac_ena~2 (
	.dataa(!col_int),
	.datab(!\Selector6~1_combout ),
	.datac(!\Selector6~2_combout ),
	.datad(!\Selector6~5_combout ),
	.datae(!\Selector7~4_combout ),
	.dataf(!\mac_ena~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mac_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mac_ena~2 .extended_lut = "off";
defparam \mac_ena~2 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \mac_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \mac_ena~3 (
	.dataa(!dreg_1),
	.datab(!Selector32),
	.datac(!\Selector0~7_combout ),
	.datad(!\Selector0~5_combout ),
	.datae(!\mac_ena~0_combout ),
	.dataf(!\mac_ena~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mac_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mac_ena~3 .extended_lut = "off";
defparam \mac_ena~3 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \mac_ena~3 .shared_arith = "off";

cyclonev_lcell_comb \stat_rden~0 (
	.dataa(!dreg_1),
	.datab(!\state.STM_TYP_IDLE~q ),
	.datac(!\Selector0~2_combout ),
	.datad(!\Selector0~5_combout ),
	.datae(!\always0~3_combout ),
	.dataf(!tx_stat_rden),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\stat_rden~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \stat_rden~0 .extended_lut = "off";
defparam \stat_rden~0 .lut_mask = 64'hFFFFDF8FFFFFFFFF;
defparam \stat_rden~0 .shared_arith = "off";

endmodule

module IoTOctopus_QSYS_altera_tse_lfsr_10 (
	reset,
	z_reg_9,
	z_reg_8,
	z_reg_7,
	z_reg_6,
	z_reg_5,
	z_reg_4,
	z_reg_3,
	z_reg_2,
	z_reg_1,
	z_reg_0,
	enable,
	tx_clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	z_reg_9;
output 	z_reg_8;
output 	z_reg_7;
output 	z_reg_6;
output 	z_reg_5;
output 	z_reg_4;
output 	z_reg_3;
output 	z_reg_2;
output 	z_reg_1;
output 	z_reg_0;
input 	enable;
input 	tx_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lfsr_o[15]~9_combout ;
wire \lfsr_o[15]~q ;
wire \lfsr_o~0_combout ;
wire \lfsr_o[0]~q ;
wire \lfsr_o[1]~5_combout ;
wire \lfsr_o[1]~q ;
wire \lfsr_o[2]~4_combout ;
wire \lfsr_o[2]~q ;
wire \lfsr_o[3]~q ;
wire \lfsr_o[4]~3_combout ;
wire \lfsr_o[4]~q ;
wire \lfsr_o[5]~q ;
wire \lfsr_o[6]~2_combout ;
wire \lfsr_o[6]~q ;
wire \lfsr_o[7]~q ;
wire \lfsr_o[8]~q ;
wire \lfsr_o[9]~1_combout ;
wire \lfsr_o[9]~q ;
wire \lfsr_o[10]~q ;
wire \lfsr_o[11]~q ;
wire \lfsr_o[12]~q ;
wire \lfsr_o[13]~8_combout ;
wire \lfsr_o[13]~q ;
wire \lfsr_o[14]~7_combout ;
wire \lfsr_o[14]~q ;
wire \z[14]~combout ;
wire \z_reg[14]~q ;
wire \z[11]~4_combout ;
wire \z[11]~combout ;
wire \z_reg[11]~q ;
wire \z[15]~combout ;
wire \z_reg[15]~q ;
wire \z[15]~6_combout ;
wire \z[10]~combout ;
wire \z_reg[10]~q ;
wire \z[14]~0_combout ;
wire \z[9]~1_combout ;
wire \z[9]~combout ;
wire \z~2_combout ;
wire \z[7]~3_combout ;
wire \z~5_combout ;
wire \z[13]~combout ;
wire \z_reg[13]~q ;
wire \z[8]~combout ;
wire \z[12]~combout ;
wire \z_reg[12]~q ;
wire \z[7]~combout ;
wire \z[6]~combout ;
wire \z[5]~combout ;
wire \z[4]~combout ;
wire \z[3]~combout ;
wire \z[2]~combout ;
wire \z[1]~combout ;
wire \z[0]~combout ;


dffeas \z_reg[9] (
	.clk(tx_clk),
	.d(\z[9]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_9),
	.prn(vcc));
defparam \z_reg[9] .is_wysiwyg = "true";
defparam \z_reg[9] .power_up = "low";

dffeas \z_reg[8] (
	.clk(tx_clk),
	.d(\z[8]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_8),
	.prn(vcc));
defparam \z_reg[8] .is_wysiwyg = "true";
defparam \z_reg[8] .power_up = "low";

dffeas \z_reg[7] (
	.clk(tx_clk),
	.d(\z[7]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_7),
	.prn(vcc));
defparam \z_reg[7] .is_wysiwyg = "true";
defparam \z_reg[7] .power_up = "low";

dffeas \z_reg[6] (
	.clk(tx_clk),
	.d(\z[6]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_6),
	.prn(vcc));
defparam \z_reg[6] .is_wysiwyg = "true";
defparam \z_reg[6] .power_up = "low";

dffeas \z_reg[5] (
	.clk(tx_clk),
	.d(\z[5]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_5),
	.prn(vcc));
defparam \z_reg[5] .is_wysiwyg = "true";
defparam \z_reg[5] .power_up = "low";

dffeas \z_reg[4] (
	.clk(tx_clk),
	.d(\z[4]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_4),
	.prn(vcc));
defparam \z_reg[4] .is_wysiwyg = "true";
defparam \z_reg[4] .power_up = "low";

dffeas \z_reg[3] (
	.clk(tx_clk),
	.d(\z[3]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_3),
	.prn(vcc));
defparam \z_reg[3] .is_wysiwyg = "true";
defparam \z_reg[3] .power_up = "low";

dffeas \z_reg[2] (
	.clk(tx_clk),
	.d(\z[2]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_2),
	.prn(vcc));
defparam \z_reg[2] .is_wysiwyg = "true";
defparam \z_reg[2] .power_up = "low";

dffeas \z_reg[1] (
	.clk(tx_clk),
	.d(\z[1]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_1),
	.prn(vcc));
defparam \z_reg[1] .is_wysiwyg = "true";
defparam \z_reg[1] .power_up = "low";

dffeas \z_reg[0] (
	.clk(tx_clk),
	.d(\z[0]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(z_reg_0),
	.prn(vcc));
defparam \z_reg[0] .is_wysiwyg = "true";
defparam \z_reg[0] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[15]~9 (
	.dataa(!\lfsr_o[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[15]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[15]~9 .extended_lut = "off";
defparam \lfsr_o[15]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[15]~9 .shared_arith = "off";

dffeas \lfsr_o[15] (
	.clk(tx_clk),
	.d(\lfsr_o[15]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[15]~q ),
	.prn(vcc));
defparam \lfsr_o[15] .is_wysiwyg = "true";
defparam \lfsr_o[15] .power_up = "low";

cyclonev_lcell_comb \lfsr_o~0 (
	.dataa(!\lfsr_o[3]~q ),
	.datab(!\lfsr_o[14]~q ),
	.datac(!\lfsr_o[12]~q ),
	.datad(!\lfsr_o[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o~0 .extended_lut = "off";
defparam \lfsr_o~0 .lut_mask = 64'h6996699669966996;
defparam \lfsr_o~0 .shared_arith = "off";

dffeas \lfsr_o[0] (
	.clk(tx_clk),
	.d(\lfsr_o~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[0]~q ),
	.prn(vcc));
defparam \lfsr_o[0] .is_wysiwyg = "true";
defparam \lfsr_o[0] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[1]~5 (
	.dataa(!\lfsr_o[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[1]~5 .extended_lut = "off";
defparam \lfsr_o[1]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[1]~5 .shared_arith = "off";

dffeas \lfsr_o[1] (
	.clk(tx_clk),
	.d(\lfsr_o[1]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[1]~q ),
	.prn(vcc));
defparam \lfsr_o[1] .is_wysiwyg = "true";
defparam \lfsr_o[1] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[2]~4 (
	.dataa(!\lfsr_o[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[2]~4 .extended_lut = "off";
defparam \lfsr_o[2]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[2]~4 .shared_arith = "off";

dffeas \lfsr_o[2] (
	.clk(tx_clk),
	.d(\lfsr_o[2]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[2]~q ),
	.prn(vcc));
defparam \lfsr_o[2] .is_wysiwyg = "true";
defparam \lfsr_o[2] .power_up = "low";

dffeas \lfsr_o[3] (
	.clk(tx_clk),
	.d(\lfsr_o[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[3]~q ),
	.prn(vcc));
defparam \lfsr_o[3] .is_wysiwyg = "true";
defparam \lfsr_o[3] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[4]~3 (
	.dataa(!\lfsr_o[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[4]~3 .extended_lut = "off";
defparam \lfsr_o[4]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[4]~3 .shared_arith = "off";

dffeas \lfsr_o[4] (
	.clk(tx_clk),
	.d(\lfsr_o[4]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[4]~q ),
	.prn(vcc));
defparam \lfsr_o[4] .is_wysiwyg = "true";
defparam \lfsr_o[4] .power_up = "low";

dffeas \lfsr_o[5] (
	.clk(tx_clk),
	.d(\lfsr_o[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[5]~q ),
	.prn(vcc));
defparam \lfsr_o[5] .is_wysiwyg = "true";
defparam \lfsr_o[5] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[6]~2 (
	.dataa(!\lfsr_o[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[6]~2 .extended_lut = "off";
defparam \lfsr_o[6]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[6]~2 .shared_arith = "off";

dffeas \lfsr_o[6] (
	.clk(tx_clk),
	.d(\lfsr_o[6]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[6]~q ),
	.prn(vcc));
defparam \lfsr_o[6] .is_wysiwyg = "true";
defparam \lfsr_o[6] .power_up = "low";

dffeas \lfsr_o[7] (
	.clk(tx_clk),
	.d(\lfsr_o[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[7]~q ),
	.prn(vcc));
defparam \lfsr_o[7] .is_wysiwyg = "true";
defparam \lfsr_o[7] .power_up = "low";

dffeas \lfsr_o[8] (
	.clk(tx_clk),
	.d(\lfsr_o[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[8]~q ),
	.prn(vcc));
defparam \lfsr_o[8] .is_wysiwyg = "true";
defparam \lfsr_o[8] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[9]~1 (
	.dataa(!\lfsr_o[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[9]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[9]~1 .extended_lut = "off";
defparam \lfsr_o[9]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[9]~1 .shared_arith = "off";

dffeas \lfsr_o[9] (
	.clk(tx_clk),
	.d(\lfsr_o[9]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[9]~q ),
	.prn(vcc));
defparam \lfsr_o[9] .is_wysiwyg = "true";
defparam \lfsr_o[9] .power_up = "low";

dffeas \lfsr_o[10] (
	.clk(tx_clk),
	.d(\lfsr_o[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[10]~q ),
	.prn(vcc));
defparam \lfsr_o[10] .is_wysiwyg = "true";
defparam \lfsr_o[10] .power_up = "low";

dffeas \lfsr_o[11] (
	.clk(tx_clk),
	.d(\lfsr_o[10]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[11]~q ),
	.prn(vcc));
defparam \lfsr_o[11] .is_wysiwyg = "true";
defparam \lfsr_o[11] .power_up = "low";

dffeas \lfsr_o[12] (
	.clk(tx_clk),
	.d(\lfsr_o[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[12]~q ),
	.prn(vcc));
defparam \lfsr_o[12] .is_wysiwyg = "true";
defparam \lfsr_o[12] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[13]~8 (
	.dataa(!\lfsr_o[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[13]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[13]~8 .extended_lut = "off";
defparam \lfsr_o[13]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[13]~8 .shared_arith = "off";

dffeas \lfsr_o[13] (
	.clk(tx_clk),
	.d(\lfsr_o[13]~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[13]~q ),
	.prn(vcc));
defparam \lfsr_o[13] .is_wysiwyg = "true";
defparam \lfsr_o[13] .power_up = "low";

cyclonev_lcell_comb \lfsr_o[14]~7 (
	.dataa(!\lfsr_o[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lfsr_o[14]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lfsr_o[14]~7 .extended_lut = "off";
defparam \lfsr_o[14]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lfsr_o[14]~7 .shared_arith = "off";

dffeas \lfsr_o[14] (
	.clk(tx_clk),
	.d(\lfsr_o[14]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\lfsr_o[14]~q ),
	.prn(vcc));
defparam \lfsr_o[14] .is_wysiwyg = "true";
defparam \lfsr_o[14] .power_up = "low";

cyclonev_lcell_comb \z[14] (
	.dataa(!z_reg_3),
	.datab(!z_reg_2),
	.datac(!\z[14]~0_combout ),
	.datad(!\lfsr_o[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[14] .extended_lut = "off";
defparam \z[14] .lut_mask = 64'h6996699669966996;
defparam \z[14] .shared_arith = "off";

dffeas \z_reg[14] (
	.clk(tx_clk),
	.d(\z[14]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\z_reg[14]~q ),
	.prn(vcc));
defparam \z_reg[14] .is_wysiwyg = "true";
defparam \z_reg[14] .power_up = "low";

cyclonev_lcell_comb \z[11]~4 (
	.dataa(!z_reg_7),
	.datab(!z_reg_0),
	.datac(!\z_reg[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[11]~4 .extended_lut = "off";
defparam \z[11]~4 .lut_mask = 64'h9696969696969696;
defparam \z[11]~4 .shared_arith = "off";

cyclonev_lcell_comb \z[11] (
	.dataa(!z_reg_3),
	.datab(!\z[11]~4_combout ),
	.datac(!\lfsr_o[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[11] .extended_lut = "off";
defparam \z[11] .lut_mask = 64'h9696969696969696;
defparam \z[11] .shared_arith = "off";

dffeas \z_reg[11] (
	.clk(tx_clk),
	.d(\z[11]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\z_reg[11]~q ),
	.prn(vcc));
defparam \z_reg[11] .is_wysiwyg = "true";
defparam \z_reg[11] .power_up = "low";

cyclonev_lcell_comb \z[15] (
	.dataa(!z_reg_3),
	.datab(!\lfsr_o[15]~q ),
	.datac(!\z[15]~6_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[15] .extended_lut = "off";
defparam \z[15] .lut_mask = 64'h9696969696969696;
defparam \z[15] .shared_arith = "off";

dffeas \z_reg[15] (
	.clk(tx_clk),
	.d(\z[15]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\z_reg[15]~q ),
	.prn(vcc));
defparam \z_reg[15] .is_wysiwyg = "true";
defparam \z_reg[15] .power_up = "low";

cyclonev_lcell_comb \z[15]~6 (
	.dataa(!z_reg_7),
	.datab(!z_reg_4),
	.datac(!\z_reg[11]~q ),
	.datad(!\z_reg[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[15]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[15]~6 .extended_lut = "off";
defparam \z[15]~6 .lut_mask = 64'h6996699669966996;
defparam \z[15]~6 .shared_arith = "off";

cyclonev_lcell_comb \z[10] (
	.dataa(!z_reg_6),
	.datab(!z_reg_3),
	.datac(!z_reg_2),
	.datad(!\z_reg[10]~q ),
	.datae(!\lfsr_o[10]~q ),
	.dataf(!\z[15]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[10] .extended_lut = "off";
defparam \z[10] .lut_mask = 64'h6996966996696996;
defparam \z[10] .shared_arith = "off";

dffeas \z_reg[10] (
	.clk(tx_clk),
	.d(\z[10]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\z_reg[10]~q ),
	.prn(vcc));
defparam \z_reg[10] .is_wysiwyg = "true";
defparam \z_reg[10] .power_up = "low";

cyclonev_lcell_comb \z[14]~0 (
	.dataa(!z_reg_6),
	.datab(!\z_reg[14]~q ),
	.datac(!\z_reg[10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[14]~0 .extended_lut = "off";
defparam \z[14]~0 .lut_mask = 64'h9696969696969696;
defparam \z[14]~0 .shared_arith = "off";

cyclonev_lcell_comb \z[9]~1 (
	.dataa(!z_reg_3),
	.datab(!z_reg_2),
	.datac(!z_reg_1),
	.datad(!\lfsr_o[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[9]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[9]~1 .extended_lut = "off";
defparam \z[9]~1 .lut_mask = 64'h6996699669966996;
defparam \z[9]~1 .shared_arith = "off";

cyclonev_lcell_comb \z[9] (
	.dataa(!z_reg_9),
	.datab(!z_reg_5),
	.datac(!\z[14]~0_combout ),
	.datad(!\z[9]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[9] .extended_lut = "off";
defparam \z[9] .lut_mask = 64'h6996699669966996;
defparam \z[9] .shared_arith = "off";

cyclonev_lcell_comb \z~2 (
	.dataa(!z_reg_4),
	.datab(!z_reg_1),
	.datac(!z_reg_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z~2 .extended_lut = "off";
defparam \z~2 .lut_mask = 64'h9696969696969696;
defparam \z~2 .shared_arith = "off";

cyclonev_lcell_comb \z[7]~3 (
	.dataa(!z_reg_8),
	.datab(!\z~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[7]~3 .extended_lut = "off";
defparam \z[7]~3 .lut_mask = 64'h6666666666666666;
defparam \z[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \z~5 (
	.dataa(!z_reg_5),
	.datab(!z_reg_2),
	.datac(!z_reg_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z~5 .extended_lut = "off";
defparam \z~5 .lut_mask = 64'h9696969696969696;
defparam \z~5 .shared_arith = "off";

cyclonev_lcell_comb \z[13] (
	.dataa(!z_reg_9),
	.datab(!\z_reg[13]~q ),
	.datac(!\z~5_combout ),
	.datad(!\lfsr_o[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[13] .extended_lut = "off";
defparam \z[13] .lut_mask = 64'h6996699669966996;
defparam \z[13] .shared_arith = "off";

dffeas \z_reg[13] (
	.clk(tx_clk),
	.d(\z[13]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\z_reg[13]~q ),
	.prn(vcc));
defparam \z_reg[13] .is_wysiwyg = "true";
defparam \z_reg[13] .power_up = "low";

cyclonev_lcell_comb \z[8] (
	.dataa(!z_reg_9),
	.datab(!z_reg_5),
	.datac(!z_reg_2),
	.datad(!\lfsr_o[8]~q ),
	.datae(!\z[7]~3_combout ),
	.dataf(!\z_reg[13]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[8] .extended_lut = "off";
defparam \z[8] .lut_mask = 64'h6996966996696996;
defparam \z[8] .shared_arith = "off";

cyclonev_lcell_comb \z[12] (
	.dataa(!z_reg_8),
	.datab(!\z~2_combout ),
	.datac(!\z_reg[12]~q ),
	.datad(!\lfsr_o[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[12] .extended_lut = "off";
defparam \z[12] .lut_mask = 64'h6996699669966996;
defparam \z[12] .shared_arith = "off";

dffeas \z_reg[12] (
	.clk(tx_clk),
	.d(\z[12]~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\z_reg[12]~q ),
	.prn(vcc));
defparam \z_reg[12] .is_wysiwyg = "true";
defparam \z_reg[12] .power_up = "low";

cyclonev_lcell_comb \z[7] (
	.dataa(!z_reg_7),
	.datab(!z_reg_3),
	.datac(!\z[7]~3_combout ),
	.datad(!\lfsr_o[7]~q ),
	.datae(!\z_reg[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[7] .extended_lut = "off";
defparam \z[7] .lut_mask = 64'h9669699696696996;
defparam \z[7] .shared_arith = "off";

cyclonev_lcell_comb \z[6] (
	.dataa(!z_reg_6),
	.datab(!z_reg_3),
	.datac(!z_reg_2),
	.datad(!\lfsr_o[6]~q ),
	.datae(!\z[11]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[6] .extended_lut = "off";
defparam \z[6] .lut_mask = 64'h9669699696696996;
defparam \z[6] .shared_arith = "off";

cyclonev_lcell_comb \z[5] (
	.dataa(!z_reg_6),
	.datab(!\z_reg[10]~q ),
	.datac(!\lfsr_o[5]~q ),
	.datad(!\z~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[5] .extended_lut = "off";
defparam \z[5] .lut_mask = 64'h6996699669966996;
defparam \z[5] .shared_arith = "off";

cyclonev_lcell_comb \z[4] (
	.dataa(!z_reg_9),
	.datab(!z_reg_5),
	.datac(!\z~2_combout ),
	.datad(!\lfsr_o[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[4] .extended_lut = "off";
defparam \z[4] .lut_mask = 64'h6996699669966996;
defparam \z[4] .shared_arith = "off";

cyclonev_lcell_comb \z[3] (
	.dataa(!z_reg_8),
	.datab(!\z[11]~4_combout ),
	.datac(!\lfsr_o[3]~q ),
	.datad(!\z_reg[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[3] .extended_lut = "off";
defparam \z[3] .lut_mask = 64'h6996699669966996;
defparam \z[3] .shared_arith = "off";

cyclonev_lcell_comb \z[2] (
	.dataa(!z_reg_7),
	.datab(!\z[14]~0_combout ),
	.datac(!\lfsr_o[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[2] .extended_lut = "off";
defparam \z[2] .lut_mask = 64'h9696969696969696;
defparam \z[2] .shared_arith = "off";

cyclonev_lcell_comb \z[1] (
	.dataa(!z_reg_9),
	.datab(!z_reg_6),
	.datac(!z_reg_5),
	.datad(!\z_reg[13]~q ),
	.datae(!\lfsr_o[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[1] .extended_lut = "off";
defparam \z[1] .lut_mask = 64'h9669699696696996;
defparam \z[1] .shared_arith = "off";

cyclonev_lcell_comb \z[0] (
	.dataa(!z_reg_8),
	.datab(!z_reg_5),
	.datac(!z_reg_4),
	.datad(!\z_reg[12]~q ),
	.datae(!\lfsr_o[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\z[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \z[0] .extended_lut = "off";
defparam \z[0] .lut_mask = 64'h9669699696696996;
defparam \z[0] .shared_arith = "off";

endmodule
