module FIFO_writer(input CLK, nRST, [63:0] DATA [3:0], DRDY,
                   output [63:0] WDATA, )